module sbox (
  input [7:0] in,
  output reg [7:0] out
);

reg [7:0] sb_mem [0:255];

always @(*) out <= sb_mem[in];


initial begin
sb_mem[8'h00] <= 8'h63;
sb_mem[8'h01] <= 8'h7c;
sb_mem[8'h02] <= 8'h77;
sb_mem[8'h03] <= 8'h7b;
sb_mem[8'h04] <= 8'hf2;
sb_mem[8'h05] <= 8'h6b;
sb_mem[8'h06] <= 8'h6f;
sb_mem[8'h07] <= 8'hc5;
sb_mem[8'h08] <= 8'h30;
sb_mem[8'h09] <= 8'h01;
sb_mem[8'h0a] <= 8'h67;
sb_mem[8'h0b] <= 8'h2b;
sb_mem[8'h0c] <= 8'hfe;
sb_mem[8'h0d] <= 8'hd7;
sb_mem[8'h0e] <= 8'hab;
sb_mem[8'h0f] <= 8'h76;
sb_mem[8'h10] <= 8'hca;
sb_mem[8'h11] <= 8'h82;
sb_mem[8'h12] <= 8'hc9;
sb_mem[8'h13] <= 8'h7d;
sb_mem[8'h14] <= 8'hfa;
sb_mem[8'h15] <= 8'h59;
sb_mem[8'h16] <= 8'h47;
sb_mem[8'h17] <= 8'hf0;
sb_mem[8'h18] <= 8'had;
sb_mem[8'h19] <= 8'hd4;
sb_mem[8'h1a] <= 8'ha2;
sb_mem[8'h1b] <= 8'haf;
sb_mem[8'h1c] <= 8'h9c;
sb_mem[8'h1d] <= 8'ha4;
sb_mem[8'h1e] <= 8'h72;
sb_mem[8'h1f] <= 8'hc0;
sb_mem[8'h20] <= 8'hb7;
sb_mem[8'h21] <= 8'hfd;
sb_mem[8'h22] <= 8'h93;
sb_mem[8'h23] <= 8'h26;
sb_mem[8'h24] <= 8'h36;
sb_mem[8'h25] <= 8'h3f;
sb_mem[8'h26] <= 8'hf7;
sb_mem[8'h27] <= 8'hcc;
sb_mem[8'h28] <= 8'h34;
sb_mem[8'h29] <= 8'ha5;
sb_mem[8'h2a] <= 8'he5;
sb_mem[8'h2b] <= 8'hf1;
sb_mem[8'h2c] <= 8'h71;
sb_mem[8'h2d] <= 8'hd8;
sb_mem[8'h2e] <= 8'h31;
sb_mem[8'h2f] <= 8'h15;
sb_mem[8'h30] <= 8'h04;
sb_mem[8'h31] <= 8'hc7;
sb_mem[8'h32] <= 8'h23;
sb_mem[8'h33] <= 8'hc3;
sb_mem[8'h34] <= 8'h18;
sb_mem[8'h35] <= 8'h96;
sb_mem[8'h36] <= 8'h05;
sb_mem[8'h37] <= 8'h9a;
sb_mem[8'h38] <= 8'h07;
sb_mem[8'h39] <= 8'h12;
sb_mem[8'h3a] <= 8'h80;
sb_mem[8'h3b] <= 8'he2;
sb_mem[8'h3c] <= 8'heb;
sb_mem[8'h3d] <= 8'h27;
sb_mem[8'h3e] <= 8'hb2;
sb_mem[8'h3f] <= 8'h75;
sb_mem[8'h40] <= 8'h09;
sb_mem[8'h41] <= 8'h83;
sb_mem[8'h42] <= 8'h2c;
sb_mem[8'h43] <= 8'h1a;
sb_mem[8'h44] <= 8'h1b;
sb_mem[8'h45] <= 8'h6e;
sb_mem[8'h46] <= 8'h5a;
sb_mem[8'h47] <= 8'ha0;
sb_mem[8'h48] <= 8'h52;
sb_mem[8'h49] <= 8'h3b;
sb_mem[8'h4a] <= 8'hd6;
sb_mem[8'h4b] <= 8'hb3;
sb_mem[8'h4c] <= 8'h29;
sb_mem[8'h4d] <= 8'he3;
sb_mem[8'h4e] <= 8'h2f;
sb_mem[8'h4f] <= 8'h84;
sb_mem[8'h50] <= 8'h53;
sb_mem[8'h51] <= 8'hd1;
sb_mem[8'h52] <= 8'h00;
sb_mem[8'h53] <= 8'hed;
sb_mem[8'h54] <= 8'h20;
sb_mem[8'h55] <= 8'hfc;
sb_mem[8'h56] <= 8'hb1;
sb_mem[8'h57] <= 8'h5b;
sb_mem[8'h58] <= 8'h6a;
sb_mem[8'h59] <= 8'hcb;
sb_mem[8'h5a] <= 8'hbe;
sb_mem[8'h5b] <= 8'h39;
sb_mem[8'h5c] <= 8'h4a;
sb_mem[8'h5d] <= 8'h4c;
sb_mem[8'h5e] <= 8'h58;
sb_mem[8'h5f] <= 8'hcf;
sb_mem[8'h60] <= 8'hd0;
sb_mem[8'h61] <= 8'hef;
sb_mem[8'h62] <= 8'haa;
sb_mem[8'h63] <= 8'hfb;
sb_mem[8'h64] <= 8'h43;
sb_mem[8'h65] <= 8'h4d;
sb_mem[8'h66] <= 8'h33;
sb_mem[8'h67] <= 8'h85;
sb_mem[8'h68] <= 8'h45;
sb_mem[8'h69] <= 8'hf9;
sb_mem[8'h6a] <= 8'h02;
sb_mem[8'h6b] <= 8'h7f;
sb_mem[8'h6c] <= 8'h50;
sb_mem[8'h6d] <= 8'h3c;
sb_mem[8'h6e] <= 8'h9f;
sb_mem[8'h6f] <= 8'ha8;
sb_mem[8'h70] <= 8'h51;
sb_mem[8'h71] <= 8'ha3;
sb_mem[8'h72] <= 8'h40;
sb_mem[8'h73] <= 8'h8f;
sb_mem[8'h74] <= 8'h92;
sb_mem[8'h75] <= 8'h9d;
sb_mem[8'h76] <= 8'h38;
sb_mem[8'h77] <= 8'hf5;
sb_mem[8'h78] <= 8'hbc;
sb_mem[8'h79] <= 8'hb6;
sb_mem[8'h7a] <= 8'hda;
sb_mem[8'h7b] <= 8'h21;
sb_mem[8'h7c] <= 8'h10;
sb_mem[8'h7d] <= 8'hff;
sb_mem[8'h7e] <= 8'hf3;
sb_mem[8'h7f] <= 8'hd2;
sb_mem[8'h80] <= 8'hcd;
sb_mem[8'h81] <= 8'h0c;
sb_mem[8'h82] <= 8'h13;
sb_mem[8'h83] <= 8'hec;
sb_mem[8'h84] <= 8'h5f;
sb_mem[8'h85] <= 8'h97;
sb_mem[8'h86] <= 8'h44;
sb_mem[8'h87] <= 8'h17;
sb_mem[8'h88] <= 8'hc4;
sb_mem[8'h89] <= 8'ha7;
sb_mem[8'h8a] <= 8'h7e;
sb_mem[8'h8b] <= 8'h3d;
sb_mem[8'h8c] <= 8'h64;
sb_mem[8'h8d] <= 8'h5d;
sb_mem[8'h8e] <= 8'h19;
sb_mem[8'h8f] <= 8'h73;
sb_mem[8'h90] <= 8'h60;
sb_mem[8'h91] <= 8'h81;
sb_mem[8'h92] <= 8'h4f;
sb_mem[8'h93] <= 8'hdc;
sb_mem[8'h94] <= 8'h22;
sb_mem[8'h95] <= 8'h2a;
sb_mem[8'h96] <= 8'h90;
sb_mem[8'h97] <= 8'h88;
sb_mem[8'h98] <= 8'h46;
sb_mem[8'h99] <= 8'hee;
sb_mem[8'h9a] <= 8'hb8;
sb_mem[8'h9b] <= 8'h14;
sb_mem[8'h9c] <= 8'hde;
sb_mem[8'h9d] <= 8'h5e;
sb_mem[8'h9e] <= 8'h0b;
sb_mem[8'h9f] <= 8'hdb;
sb_mem[8'ha0] <= 8'he0;
sb_mem[8'ha1] <= 8'h32;
sb_mem[8'ha2] <= 8'h3a;
sb_mem[8'ha3] <= 8'h0a;
sb_mem[8'ha4] <= 8'h49;
sb_mem[8'ha5] <= 8'h06;
sb_mem[8'ha6] <= 8'h24;
sb_mem[8'ha7] <= 8'h5c;
sb_mem[8'ha8] <= 8'hc2;
sb_mem[8'ha9] <= 8'hd3;
sb_mem[8'haa] <= 8'hac;
sb_mem[8'hab] <= 8'h62;
sb_mem[8'hac] <= 8'h91;
sb_mem[8'had] <= 8'h95;
sb_mem[8'hae] <= 8'he4;
sb_mem[8'haf] <= 8'h79;
sb_mem[8'hb0] <= 8'he7;
sb_mem[8'hb1] <= 8'hc8;
sb_mem[8'hb2] <= 8'h37;
sb_mem[8'hb3] <= 8'h6d;
sb_mem[8'hb4] <= 8'h8d;
sb_mem[8'hb5] <= 8'hd5;
sb_mem[8'hb6] <= 8'h4e;
sb_mem[8'hb7] <= 8'ha9;
sb_mem[8'hb8] <= 8'h6c;
sb_mem[8'hb9] <= 8'h56;
sb_mem[8'hba] <= 8'hf4;
sb_mem[8'hbb] <= 8'hea;
sb_mem[8'hbc] <= 8'h65;
sb_mem[8'hbd] <= 8'h7a;
sb_mem[8'hbe] <= 8'hae;
sb_mem[8'hbf] <= 8'h08;
sb_mem[8'hc0] <= 8'hba;
sb_mem[8'hc1] <= 8'h78;
sb_mem[8'hc2] <= 8'h25;
sb_mem[8'hc3] <= 8'h2e;
sb_mem[8'hc4] <= 8'h1c;
sb_mem[8'hc5] <= 8'ha6;
sb_mem[8'hc6] <= 8'hb4;
sb_mem[8'hc7] <= 8'hc6;
sb_mem[8'hc8] <= 8'he8;
sb_mem[8'hc9] <= 8'hdd;
sb_mem[8'hca] <= 8'h74;
sb_mem[8'hcb] <= 8'h1f;
sb_mem[8'hcc] <= 8'h4b;
sb_mem[8'hcd] <= 8'hbd;
sb_mem[8'hce] <= 8'h8b;
sb_mem[8'hcf] <= 8'h8a;
sb_mem[8'hd0] <= 8'h70;
sb_mem[8'hd1] <= 8'h3e;
sb_mem[8'hd2] <= 8'hb5;
sb_mem[8'hd3] <= 8'h66;
sb_mem[8'hd4] <= 8'h48;
sb_mem[8'hd5] <= 8'h03;
sb_mem[8'hd6] <= 8'hf6;
sb_mem[8'hd7] <= 8'h0e;
sb_mem[8'hd8] <= 8'h61;
sb_mem[8'hd9] <= 8'h35;
sb_mem[8'hda] <= 8'h57;
sb_mem[8'hdb] <= 8'hb9;
sb_mem[8'hdc] <= 8'h86;
sb_mem[8'hdd] <= 8'hc1;
sb_mem[8'hde] <= 8'h1d;
sb_mem[8'hdf] <= 8'h9e;
sb_mem[8'he0] <= 8'he1;
sb_mem[8'he1] <= 8'hf8;
sb_mem[8'he2] <= 8'h98;
sb_mem[8'he3] <= 8'h11;
sb_mem[8'he4] <= 8'h69;
sb_mem[8'he5] <= 8'hd9;
sb_mem[8'he6] <= 8'h8e;
sb_mem[8'he7] <= 8'h94;
sb_mem[8'he8] <= 8'h9b;
sb_mem[8'he9] <= 8'h1e;
sb_mem[8'hea] <= 8'h87;
sb_mem[8'heb] <= 8'he9;
sb_mem[8'hec] <= 8'hce;
sb_mem[8'hed] <= 8'h55;
sb_mem[8'hee] <= 8'h28;
sb_mem[8'hef] <= 8'hdf;
sb_mem[8'hf0] <= 8'h8c;
sb_mem[8'hf1] <= 8'ha1;
sb_mem[8'hf2] <= 8'h89;
sb_mem[8'hf3] <= 8'h0d;
sb_mem[8'hf4] <= 8'hbf;
sb_mem[8'hf5] <= 8'he6;
sb_mem[8'hf6] <= 8'h42;
sb_mem[8'hf7] <= 8'h68;
sb_mem[8'hf8] <= 8'h41;
sb_mem[8'hf9] <= 8'h99;
sb_mem[8'hfa] <= 8'h2d;
sb_mem[8'hfb] <= 8'h0f;
sb_mem[8'hfc] <= 8'hb0;
sb_mem[8'hfd] <= 8'h54;
sb_mem[8'hfe] <= 8'hbb;
sb_mem[8'hff] <= 8'h16;
end



endmodule 
