module M13 (
  input [7:0] in,
  output reg [7:0] out
);

reg [7:0] m13_mem [0:255];

always @(*) out = m13_mem[in];

initial begin
m13_mem[8'h00] <= 8'h00;
m13_mem[8'h01] <= 8'h0d;
m13_mem[8'h02] <= 8'h1a;
m13_mem[8'h03] <= 8'h17;
m13_mem[8'h04] <= 8'h34;
m13_mem[8'h05] <= 8'h39;
m13_mem[8'h06] <= 8'h2e;
m13_mem[8'h07] <= 8'h23;
m13_mem[8'h08] <= 8'h68;
m13_mem[8'h09] <= 8'h65;
m13_mem[8'h0a] <= 8'h72;
m13_mem[8'h0b] <= 8'h7f;
m13_mem[8'h0c] <= 8'h5c;
m13_mem[8'h0d] <= 8'h51;
m13_mem[8'h0e] <= 8'h46;
m13_mem[8'h0f] <= 8'h4b;
m13_mem[8'h10] <= 8'hd0;
m13_mem[8'h11] <= 8'hdd;
m13_mem[8'h12] <= 8'hca;
m13_mem[8'h13] <= 8'hc7;
m13_mem[8'h14] <= 8'he4;
m13_mem[8'h15] <= 8'he9;
m13_mem[8'h16] <= 8'hfe;
m13_mem[8'h17] <= 8'hf3;
m13_mem[8'h18] <= 8'hb8;
m13_mem[8'h19] <= 8'hb5;
m13_mem[8'h1a] <= 8'ha2;
m13_mem[8'h1b] <= 8'haf;
m13_mem[8'h1c] <= 8'h8c;
m13_mem[8'h1d] <= 8'h81;
m13_mem[8'h1e] <= 8'h96;
m13_mem[8'h1f] <= 8'h9b;
m13_mem[8'h20] <= 8'hbb;
m13_mem[8'h21] <= 8'hb6;
m13_mem[8'h22] <= 8'ha1;
m13_mem[8'h23] <= 8'hac;
m13_mem[8'h24] <= 8'h8f;
m13_mem[8'h25] <= 8'h82;
m13_mem[8'h26] <= 8'h95;
m13_mem[8'h27] <= 8'h98;
m13_mem[8'h28] <= 8'hd3;
m13_mem[8'h29] <= 8'hde;
m13_mem[8'h2a] <= 8'hc9;
m13_mem[8'h2b] <= 8'hc4;
m13_mem[8'h2c] <= 8'he7;
m13_mem[8'h2d] <= 8'hea;
m13_mem[8'h2e] <= 8'hfd;
m13_mem[8'h2f] <= 8'hf0;
m13_mem[8'h30] <= 8'h6b;
m13_mem[8'h31] <= 8'h66;
m13_mem[8'h32] <= 8'h71;
m13_mem[8'h33] <= 8'h7c;
m13_mem[8'h34] <= 8'h5f;
m13_mem[8'h35] <= 8'h52;
m13_mem[8'h36] <= 8'h45;
m13_mem[8'h37] <= 8'h48;
m13_mem[8'h38] <= 8'h03;
m13_mem[8'h39] <= 8'h0e;
m13_mem[8'h3a] <= 8'h19;
m13_mem[8'h3b] <= 8'h14;
m13_mem[8'h3c] <= 8'h37;
m13_mem[8'h3d] <= 8'h3a;
m13_mem[8'h3e] <= 8'h2d;
m13_mem[8'h3f] <= 8'h20;
m13_mem[8'h40] <= 8'h6d;
m13_mem[8'h41] <= 8'h60;
m13_mem[8'h42] <= 8'h77;
m13_mem[8'h43] <= 8'h7a;
m13_mem[8'h44] <= 8'h59;
m13_mem[8'h45] <= 8'h54;
m13_mem[8'h46] <= 8'h43;
m13_mem[8'h47] <= 8'h4e;
m13_mem[8'h48] <= 8'h05;
m13_mem[8'h49] <= 8'h08;
m13_mem[8'h4a] <= 8'h1f;
m13_mem[8'h4b] <= 8'h12;
m13_mem[8'h4c] <= 8'h31;
m13_mem[8'h4d] <= 8'h3c;
m13_mem[8'h4e] <= 8'h2b;
m13_mem[8'h4f] <= 8'h26;
m13_mem[8'h50] <= 8'hbd;
m13_mem[8'h51] <= 8'hb0;
m13_mem[8'h52] <= 8'ha7;
m13_mem[8'h53] <= 8'haa;
m13_mem[8'h54] <= 8'h89;
m13_mem[8'h55] <= 8'h84;
m13_mem[8'h56] <= 8'h93;
m13_mem[8'h57] <= 8'h9e;
m13_mem[8'h58] <= 8'hd5;
m13_mem[8'h59] <= 8'hd8;
m13_mem[8'h5a] <= 8'hcf;
m13_mem[8'h5b] <= 8'hc2;
m13_mem[8'h5c] <= 8'he1;
m13_mem[8'h5d] <= 8'hec;
m13_mem[8'h5e] <= 8'hfb;
m13_mem[8'h5f] <= 8'hf6;
m13_mem[8'h60] <= 8'hd6;
m13_mem[8'h61] <= 8'hdb;
m13_mem[8'h62] <= 8'hcc;
m13_mem[8'h63] <= 8'hc1;
m13_mem[8'h64] <= 8'he2;
m13_mem[8'h65] <= 8'hef;
m13_mem[8'h66] <= 8'hf8;
m13_mem[8'h67] <= 8'hf5;
m13_mem[8'h68] <= 8'hbe;
m13_mem[8'h69] <= 8'hb3;
m13_mem[8'h6a] <= 8'ha4;
m13_mem[8'h6b] <= 8'ha9;
m13_mem[8'h6c] <= 8'h8a;
m13_mem[8'h6d] <= 8'h87;
m13_mem[8'h6e] <= 8'h90;
m13_mem[8'h6f] <= 8'h9d;
m13_mem[8'h70] <= 8'h06;
m13_mem[8'h71] <= 8'h0b;
m13_mem[8'h72] <= 8'h1c;
m13_mem[8'h73] <= 8'h11;
m13_mem[8'h74] <= 8'h32;
m13_mem[8'h75] <= 8'h3f;
m13_mem[8'h76] <= 8'h28;
m13_mem[8'h77] <= 8'h25;
m13_mem[8'h78] <= 8'h6e;
m13_mem[8'h79] <= 8'h63;
m13_mem[8'h7a] <= 8'h74;
m13_mem[8'h7b] <= 8'h79;
m13_mem[8'h7c] <= 8'h5a;
m13_mem[8'h7d] <= 8'h57;
m13_mem[8'h7e] <= 8'h40;
m13_mem[8'h7f] <= 8'h4d;
m13_mem[8'h80] <= 8'hda;
m13_mem[8'h81] <= 8'hd7;
m13_mem[8'h82] <= 8'hc0;
m13_mem[8'h83] <= 8'hcd;
m13_mem[8'h84] <= 8'hee;
m13_mem[8'h85] <= 8'he3;
m13_mem[8'h86] <= 8'hf4;
m13_mem[8'h87] <= 8'hf9;
m13_mem[8'h88] <= 8'hb2;
m13_mem[8'h89] <= 8'hbf;
m13_mem[8'h8a] <= 8'ha8;
m13_mem[8'h8b] <= 8'ha5;
m13_mem[8'h8c] <= 8'h86;
m13_mem[8'h8d] <= 8'h8b;
m13_mem[8'h8e] <= 8'h9c;
m13_mem[8'h8f] <= 8'h91;
m13_mem[8'h90] <= 8'h0a;
m13_mem[8'h91] <= 8'h07;
m13_mem[8'h92] <= 8'h10;
m13_mem[8'h93] <= 8'h1d;
m13_mem[8'h94] <= 8'h3e;
m13_mem[8'h95] <= 8'h33;
m13_mem[8'h96] <= 8'h24;
m13_mem[8'h97] <= 8'h29;
m13_mem[8'h98] <= 8'h62;
m13_mem[8'h99] <= 8'h6f;
m13_mem[8'h9a] <= 8'h78;
m13_mem[8'h9b] <= 8'h75;
m13_mem[8'h9c] <= 8'h56;
m13_mem[8'h9d] <= 8'h5b;
m13_mem[8'h9e] <= 8'h4c;
m13_mem[8'h9f] <= 8'h41;
m13_mem[8'ha0] <= 8'h61;
m13_mem[8'ha1] <= 8'h6c;
m13_mem[8'ha2] <= 8'h7b;
m13_mem[8'ha3] <= 8'h76;
m13_mem[8'ha4] <= 8'h55;
m13_mem[8'ha5] <= 8'h58;
m13_mem[8'ha6] <= 8'h4f;
m13_mem[8'ha7] <= 8'h42;
m13_mem[8'ha8] <= 8'h09;
m13_mem[8'ha9] <= 8'h04;
m13_mem[8'haa] <= 8'h13;
m13_mem[8'hab] <= 8'h1e;
m13_mem[8'hac] <= 8'h3d;
m13_mem[8'had] <= 8'h30;
m13_mem[8'hae] <= 8'h27;
m13_mem[8'haf] <= 8'h2a;
m13_mem[8'hb0] <= 8'hb1;
m13_mem[8'hb1] <= 8'hbc;
m13_mem[8'hb2] <= 8'hab;
m13_mem[8'hb3] <= 8'ha6;
m13_mem[8'hb4] <= 8'h85;
m13_mem[8'hb5] <= 8'h88;
m13_mem[8'hb6] <= 8'h9f;
m13_mem[8'hb7] <= 8'h92;
m13_mem[8'hb8] <= 8'hd9;
m13_mem[8'hb9] <= 8'hd4;
m13_mem[8'hba] <= 8'hc3;
m13_mem[8'hbb] <= 8'hce;
m13_mem[8'hbc] <= 8'hed;
m13_mem[8'hbd] <= 8'he0;
m13_mem[8'hbe] <= 8'hf7;
m13_mem[8'hbf] <= 8'hfa;
m13_mem[8'hc0] <= 8'hb7;
m13_mem[8'hc1] <= 8'hba;
m13_mem[8'hc2] <= 8'had;
m13_mem[8'hc3] <= 8'ha0;
m13_mem[8'hc4] <= 8'h83;
m13_mem[8'hc5] <= 8'h8e;
m13_mem[8'hc6] <= 8'h99;
m13_mem[8'hc7] <= 8'h94;
m13_mem[8'hc8] <= 8'hdf;
m13_mem[8'hc9] <= 8'hd2;
m13_mem[8'hca] <= 8'hc5;
m13_mem[8'hcb] <= 8'hc8;
m13_mem[8'hcc] <= 8'heb;
m13_mem[8'hcd] <= 8'he6;
m13_mem[8'hce] <= 8'hf1;
m13_mem[8'hcf] <= 8'hfc;
m13_mem[8'hd0] <= 8'h67;
m13_mem[8'hd1] <= 8'h6a;
m13_mem[8'hd2] <= 8'h7d;
m13_mem[8'hd3] <= 8'h70;
m13_mem[8'hd4] <= 8'h53;
m13_mem[8'hd5] <= 8'h5e;
m13_mem[8'hd6] <= 8'h49;
m13_mem[8'hd7] <= 8'h44;
m13_mem[8'hd8] <= 8'h0f;
m13_mem[8'hd9] <= 8'h02;
m13_mem[8'hda] <= 8'h15;
m13_mem[8'hdb] <= 8'h18;
m13_mem[8'hdc] <= 8'h3b;
m13_mem[8'hdd] <= 8'h36;
m13_mem[8'hde] <= 8'h21;
m13_mem[8'hdf] <= 8'h2c;
m13_mem[8'he0] <= 8'h0c;
m13_mem[8'he1] <= 8'h01;
m13_mem[8'he2] <= 8'h16;
m13_mem[8'he3] <= 8'h1b;
m13_mem[8'he4] <= 8'h38;
m13_mem[8'he5] <= 8'h35;
m13_mem[8'he6] <= 8'h22;
m13_mem[8'he7] <= 8'h2f;
m13_mem[8'he8] <= 8'h64;
m13_mem[8'he9] <= 8'h69;
m13_mem[8'hea] <= 8'h7e;
m13_mem[8'heb] <= 8'h73;
m13_mem[8'hec] <= 8'h50;
m13_mem[8'hed] <= 8'h5d;
m13_mem[8'hee] <= 8'h4a;
m13_mem[8'hef] <= 8'h47;
m13_mem[8'hf0] <= 8'hdc;
m13_mem[8'hf1] <= 8'hd1;
m13_mem[8'hf2] <= 8'hc6;
m13_mem[8'hf3] <= 8'hcb;
m13_mem[8'hf4] <= 8'he8;
m13_mem[8'hf5] <= 8'he5;
m13_mem[8'hf6] <= 8'hf2;
m13_mem[8'hf7] <= 8'hff;
m13_mem[8'hf8] <= 8'hb4;
m13_mem[8'hf9] <= 8'hb9;
m13_mem[8'hfa] <= 8'hae;
m13_mem[8'hfb] <= 8'ha3;
m13_mem[8'hfc] <= 8'h80;
m13_mem[8'hfd] <= 8'h8d;
m13_mem[8'hfe] <= 8'h9a;
m13_mem[8'hff] <= 8'h97;
end  


endmodule
