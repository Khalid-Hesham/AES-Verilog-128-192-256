module M3 (
  input [7:0] in,
  output reg [7:0] out
);

reg [7:0] m3_mem [0:255] ;

always @(*) out = m3_mem[in];


initial begin
m3_mem[8'h00] <= 8'h00;
m3_mem[8'h01] <= 8'h03;
m3_mem[8'h02] <= 8'h06;
m3_mem[8'h03] <= 8'h05;
m3_mem[8'h04] <= 8'h0c;
m3_mem[8'h05] <= 8'h0f;
m3_mem[8'h06] <= 8'h0a;
m3_mem[8'h07] <= 8'h09;
m3_mem[8'h08] <= 8'h18;
m3_mem[8'h09] <= 8'h1b;
m3_mem[8'h0a] <= 8'h1e;
m3_mem[8'h0b] <= 8'h1d;
m3_mem[8'h0c] <= 8'h14;
m3_mem[8'h0d] <= 8'h17;
m3_mem[8'h0e] <= 8'h12;
m3_mem[8'h0f] <= 8'h11;
m3_mem[8'h10] <= 8'h30;
m3_mem[8'h11] <= 8'h33;
m3_mem[8'h12] <= 8'h36;
m3_mem[8'h13] <= 8'h35;
m3_mem[8'h14] <= 8'h3c;
m3_mem[8'h15] <= 8'h3f;
m3_mem[8'h16] <= 8'h3a;
m3_mem[8'h17] <= 8'h39;
m3_mem[8'h18] <= 8'h28;
m3_mem[8'h19] <= 8'h2b;
m3_mem[8'h1a] <= 8'h2e;
m3_mem[8'h1b] <= 8'h2d;
m3_mem[8'h1c] <= 8'h24;
m3_mem[8'h1d] <= 8'h27;
m3_mem[8'h1e] <= 8'h22;
m3_mem[8'h1f] <= 8'h21;
m3_mem[8'h20] <= 8'h60;
m3_mem[8'h21] <= 8'h63;
m3_mem[8'h22] <= 8'h66;
m3_mem[8'h23] <= 8'h65;
m3_mem[8'h24] <= 8'h6c;
m3_mem[8'h25] <= 8'h6f;
m3_mem[8'h26] <= 8'h6a;
m3_mem[8'h27] <= 8'h69;
m3_mem[8'h28] <= 8'h78;
m3_mem[8'h29] <= 8'h7b;
m3_mem[8'h2a] <= 8'h7e;
m3_mem[8'h2b] <= 8'h7d;
m3_mem[8'h2c] <= 8'h74;
m3_mem[8'h2d] <= 8'h77;
m3_mem[8'h2e] <= 8'h72;
m3_mem[8'h2f] <= 8'h71;
m3_mem[8'h30] <= 8'h50;
m3_mem[8'h31] <= 8'h53;
m3_mem[8'h32] <= 8'h56;
m3_mem[8'h33] <= 8'h55;
m3_mem[8'h34] <= 8'h5c;
m3_mem[8'h35] <= 8'h5f;
m3_mem[8'h36] <= 8'h5a;
m3_mem[8'h37] <= 8'h59;
m3_mem[8'h38] <= 8'h48;
m3_mem[8'h39] <= 8'h4b;
m3_mem[8'h3a] <= 8'h4e;
m3_mem[8'h3b] <= 8'h4d;
m3_mem[8'h3c] <= 8'h44;
m3_mem[8'h3d] <= 8'h47;
m3_mem[8'h3e] <= 8'h42;
m3_mem[8'h3f] <= 8'h41;
m3_mem[8'h40] <= 8'hc0;
m3_mem[8'h41] <= 8'hc3;
m3_mem[8'h42] <= 8'hc6;
m3_mem[8'h43] <= 8'hc5;
m3_mem[8'h44] <= 8'hcc;
m3_mem[8'h45] <= 8'hcf;
m3_mem[8'h46] <= 8'hca;
m3_mem[8'h47] <= 8'hc9;
m3_mem[8'h48] <= 8'hd8;
m3_mem[8'h49] <= 8'hdb;
m3_mem[8'h4a] <= 8'hde;
m3_mem[8'h4b] <= 8'hdd;
m3_mem[8'h4c] <= 8'hd4;
m3_mem[8'h4d] <= 8'hd7;
m3_mem[8'h4e] <= 8'hd2;
m3_mem[8'h4f] <= 8'hd1;
m3_mem[8'h50] <= 8'hf0;
m3_mem[8'h51] <= 8'hf3;
m3_mem[8'h52] <= 8'hf6;
m3_mem[8'h53] <= 8'hf5;
m3_mem[8'h54] <= 8'hfc;
m3_mem[8'h55] <= 8'hff;
m3_mem[8'h56] <= 8'hfa;
m3_mem[8'h57] <= 8'hf9;
m3_mem[8'h58] <= 8'he8;
m3_mem[8'h59] <= 8'heb;
m3_mem[8'h5a] <= 8'hee;
m3_mem[8'h5b] <= 8'hed;
m3_mem[8'h5c] <= 8'he4;
m3_mem[8'h5d] <= 8'he7;
m3_mem[8'h5e] <= 8'he2;
m3_mem[8'h5f] <= 8'he1;
m3_mem[8'h60] <= 8'ha0;
m3_mem[8'h61] <= 8'ha3;
m3_mem[8'h62] <= 8'ha6;
m3_mem[8'h63] <= 8'ha5;
m3_mem[8'h64] <= 8'hac;
m3_mem[8'h65] <= 8'haf;
m3_mem[8'h66] <= 8'haa;
m3_mem[8'h67] <= 8'ha9;
m3_mem[8'h68] <= 8'hb8;
m3_mem[8'h69] <= 8'hbb;
m3_mem[8'h6a] <= 8'hbe;
m3_mem[8'h6b] <= 8'hbd;
m3_mem[8'h6c] <= 8'hb4;
m3_mem[8'h6d] <= 8'hb7;
m3_mem[8'h6e] <= 8'hb2;
m3_mem[8'h6f] <= 8'hb1;
m3_mem[8'h70] <= 8'h90;
m3_mem[8'h71] <= 8'h93;
m3_mem[8'h72] <= 8'h96;
m3_mem[8'h73] <= 8'h95;
m3_mem[8'h74] <= 8'h9c;
m3_mem[8'h75] <= 8'h9f;
m3_mem[8'h76] <= 8'h9a;
m3_mem[8'h77] <= 8'h99;
m3_mem[8'h78] <= 8'h88;
m3_mem[8'h79] <= 8'h8b;
m3_mem[8'h7a] <= 8'h8e;
m3_mem[8'h7b] <= 8'h8d;
m3_mem[8'h7c] <= 8'h84;
m3_mem[8'h7d] <= 8'h87;
m3_mem[8'h7e] <= 8'h82;
m3_mem[8'h7f] <= 8'h81;
m3_mem[8'h80] <= 8'h9b;
m3_mem[8'h81] <= 8'h98;
m3_mem[8'h82] <= 8'h9d;
m3_mem[8'h83] <= 8'h9e;
m3_mem[8'h84] <= 8'h97;
m3_mem[8'h85] <= 8'h94;
m3_mem[8'h86] <= 8'h91;
m3_mem[8'h87] <= 8'h92;
m3_mem[8'h88] <= 8'h83;
m3_mem[8'h89] <= 8'h80;
m3_mem[8'h8a] <= 8'h85;
m3_mem[8'h8b] <= 8'h86;
m3_mem[8'h8c] <= 8'h8f;
m3_mem[8'h8d] <= 8'h8c;
m3_mem[8'h8e] <= 8'h89;
m3_mem[8'h8f] <= 8'h8a;
m3_mem[8'h90] <= 8'hab;
m3_mem[8'h91] <= 8'ha8;
m3_mem[8'h92] <= 8'had;
m3_mem[8'h93] <= 8'hae;
m3_mem[8'h94] <= 8'ha7;
m3_mem[8'h95] <= 8'ha4;
m3_mem[8'h96] <= 8'ha1;
m3_mem[8'h97] <= 8'ha2;
m3_mem[8'h98] <= 8'hb3;
m3_mem[8'h99] <= 8'hb0;
m3_mem[8'h9a] <= 8'hb5;
m3_mem[8'h9b] <= 8'hb6;
m3_mem[8'h9c] <= 8'hbf;
m3_mem[8'h9d] <= 8'hbc;
m3_mem[8'h9e] <= 8'hb9;
m3_mem[8'h9f] <= 8'hba;
m3_mem[8'ha0] <= 8'hfb;
m3_mem[8'ha1] <= 8'hf8;
m3_mem[8'ha2] <= 8'hfd;
m3_mem[8'ha3] <= 8'hfe;
m3_mem[8'ha4] <= 8'hf7;
m3_mem[8'ha5] <= 8'hf4;
m3_mem[8'ha6] <= 8'hf1;
m3_mem[8'ha7] <= 8'hf2;
m3_mem[8'ha8] <= 8'he3;
m3_mem[8'ha9] <= 8'he0;
m3_mem[8'haa] <= 8'he5;
m3_mem[8'hab] <= 8'he6;
m3_mem[8'hac] <= 8'hef;
m3_mem[8'had] <= 8'hec;
m3_mem[8'hae] <= 8'he9;
m3_mem[8'haf] <= 8'hea;
m3_mem[8'hb0] <= 8'hcb;
m3_mem[8'hb1] <= 8'hc8;
m3_mem[8'hb2] <= 8'hcd;
m3_mem[8'hb3] <= 8'hce;
m3_mem[8'hb4] <= 8'hc7;
m3_mem[8'hb5] <= 8'hc4;
m3_mem[8'hb6] <= 8'hc1;
m3_mem[8'hb7] <= 8'hc2;
m3_mem[8'hb8] <= 8'hd3;
m3_mem[8'hb9] <= 8'hd0;
m3_mem[8'hba] <= 8'hd5;
m3_mem[8'hbb] <= 8'hd6;
m3_mem[8'hbc] <= 8'hdf;
m3_mem[8'hbd] <= 8'hdc;
m3_mem[8'hbe] <= 8'hd9;
m3_mem[8'hbf] <= 8'hda;
m3_mem[8'hc0] <= 8'h5b;
m3_mem[8'hc1] <= 8'h58;
m3_mem[8'hc2] <= 8'h5d;
m3_mem[8'hc3] <= 8'h5e;
m3_mem[8'hc4] <= 8'h57;
m3_mem[8'hc5] <= 8'h54;
m3_mem[8'hc6] <= 8'h51;
m3_mem[8'hc7] <= 8'h52;
m3_mem[8'hc8] <= 8'h43;
m3_mem[8'hc9] <= 8'h40;
m3_mem[8'hca] <= 8'h45;
m3_mem[8'hcb] <= 8'h46;
m3_mem[8'hcc] <= 8'h4f;
m3_mem[8'hcd] <= 8'h4c;
m3_mem[8'hce] <= 8'h49;
m3_mem[8'hcf] <= 8'h4a;
m3_mem[8'hd0] <= 8'h6b;
m3_mem[8'hd1] <= 8'h68;
m3_mem[8'hd2] <= 8'h6d;
m3_mem[8'hd3] <= 8'h6e;
m3_mem[8'hd4] <= 8'h67;
m3_mem[8'hd5] <= 8'h64;
m3_mem[8'hd6] <= 8'h61;
m3_mem[8'hd7] <= 8'h62;
m3_mem[8'hd8] <= 8'h73;
m3_mem[8'hd9] <= 8'h70;
m3_mem[8'hda] <= 8'h75;
m3_mem[8'hdb] <= 8'h76;
m3_mem[8'hdc] <= 8'h7f;
m3_mem[8'hdd] <= 8'h7c;
m3_mem[8'hde] <= 8'h79;
m3_mem[8'hdf] <= 8'h7a;
m3_mem[8'he0] <= 8'h3b;
m3_mem[8'he1] <= 8'h38;
m3_mem[8'he2] <= 8'h3d;
m3_mem[8'he3] <= 8'h3e;
m3_mem[8'he4] <= 8'h37;
m3_mem[8'he5] <= 8'h34;
m3_mem[8'he6] <= 8'h31;
m3_mem[8'he7] <= 8'h32;
m3_mem[8'he8] <= 8'h23;
m3_mem[8'he9] <= 8'h20;
m3_mem[8'hea] <= 8'h25;
m3_mem[8'heb] <= 8'h26;
m3_mem[8'hec] <= 8'h2f;
m3_mem[8'hed] <= 8'h2c;
m3_mem[8'hee] <= 8'h29;
m3_mem[8'hef] <= 8'h2a;
m3_mem[8'hf0] <= 8'h0b;
m3_mem[8'hf1] <= 8'h08;
m3_mem[8'hf2] <= 8'h0d;
m3_mem[8'hf3] <= 8'h0e;
m3_mem[8'hf4] <= 8'h07;
m3_mem[8'hf5] <= 8'h04;
m3_mem[8'hf6] <= 8'h01;
m3_mem[8'hf7] <= 8'h02;
m3_mem[8'hf8] <= 8'h13;
m3_mem[8'hf9] <= 8'h10;
m3_mem[8'hfa] <= 8'h15;
m3_mem[8'hfb] <= 8'h16;
m3_mem[8'hfc] <= 8'h1f;
m3_mem[8'hfd] <= 8'h1c;
m3_mem[8'hfe] <= 8'h19;
m3_mem[8'hff] <= 8'h1a;
end  

endmodule
