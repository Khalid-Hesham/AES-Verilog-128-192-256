module M11 (
  input [7:0] in,
  output reg [7:0] out
);

reg [7:0] m11_mem [0:255];

always @(*) out = m11_mem[in];

initial begin
m11_mem[8'h00] <= 8'h00;
m11_mem[8'h01] <= 8'h0b;
m11_mem[8'h02] <= 8'h16;
m11_mem[8'h03] <= 8'h1d;
m11_mem[8'h04] <= 8'h2c;
m11_mem[8'h05] <= 8'h27;
m11_mem[8'h06] <= 8'h3a;
m11_mem[8'h07] <= 8'h31;
m11_mem[8'h08] <= 8'h58;
m11_mem[8'h09] <= 8'h53;
m11_mem[8'h0a] <= 8'h4e;
m11_mem[8'h0b] <= 8'h45;
m11_mem[8'h0c] <= 8'h74;
m11_mem[8'h0d] <= 8'h7f;
m11_mem[8'h0e] <= 8'h62;
m11_mem[8'h0f] <= 8'h69;
m11_mem[8'h10] <= 8'hb0;
m11_mem[8'h11] <= 8'hbb;
m11_mem[8'h12] <= 8'ha6;
m11_mem[8'h13] <= 8'had;
m11_mem[8'h14] <= 8'h9c;
m11_mem[8'h15] <= 8'h97;
m11_mem[8'h16] <= 8'h8a;
m11_mem[8'h17] <= 8'h81;
m11_mem[8'h18] <= 8'he8;
m11_mem[8'h19] <= 8'he3;
m11_mem[8'h1a] <= 8'hfe;
m11_mem[8'h1b] <= 8'hf5;
m11_mem[8'h1c] <= 8'hc4;
m11_mem[8'h1d] <= 8'hcf;
m11_mem[8'h1e] <= 8'hd2;
m11_mem[8'h1f] <= 8'hd9;
m11_mem[8'h20] <= 8'h7b;
m11_mem[8'h21] <= 8'h70;
m11_mem[8'h22] <= 8'h6d;
m11_mem[8'h23] <= 8'h66;
m11_mem[8'h24] <= 8'h57;
m11_mem[8'h25] <= 8'h5c;
m11_mem[8'h26] <= 8'h41;
m11_mem[8'h27] <= 8'h4a;
m11_mem[8'h28] <= 8'h23;
m11_mem[8'h29] <= 8'h28;
m11_mem[8'h2a] <= 8'h35;
m11_mem[8'h2b] <= 8'h3e;
m11_mem[8'h2c] <= 8'h0f;
m11_mem[8'h2d] <= 8'h04;
m11_mem[8'h2e] <= 8'h19;
m11_mem[8'h2f] <= 8'h12;
m11_mem[8'h30] <= 8'hcb;
m11_mem[8'h31] <= 8'hc0;
m11_mem[8'h32] <= 8'hdd;
m11_mem[8'h33] <= 8'hd6;
m11_mem[8'h34] <= 8'he7;
m11_mem[8'h35] <= 8'hec;
m11_mem[8'h36] <= 8'hf1;
m11_mem[8'h37] <= 8'hfa;
m11_mem[8'h38] <= 8'h93;
m11_mem[8'h39] <= 8'h98;
m11_mem[8'h3a] <= 8'h85;
m11_mem[8'h3b] <= 8'h8e;
m11_mem[8'h3c] <= 8'hbf;
m11_mem[8'h3d] <= 8'hb4;
m11_mem[8'h3e] <= 8'ha9;
m11_mem[8'h3f] <= 8'ha2;
m11_mem[8'h40] <= 8'hf6;
m11_mem[8'h41] <= 8'hfd;
m11_mem[8'h42] <= 8'he0;
m11_mem[8'h43] <= 8'heb;
m11_mem[8'h44] <= 8'hda;
m11_mem[8'h45] <= 8'hd1;
m11_mem[8'h46] <= 8'hcc;
m11_mem[8'h47] <= 8'hc7;
m11_mem[8'h48] <= 8'hae;
m11_mem[8'h49] <= 8'ha5;
m11_mem[8'h4a] <= 8'hb8;
m11_mem[8'h4b] <= 8'hb3;
m11_mem[8'h4c] <= 8'h82;
m11_mem[8'h4d] <= 8'h89;
m11_mem[8'h4e] <= 8'h94;
m11_mem[8'h4f] <= 8'h9f;
m11_mem[8'h50] <= 8'h46;
m11_mem[8'h51] <= 8'h4d;
m11_mem[8'h52] <= 8'h50;
m11_mem[8'h53] <= 8'h5b;
m11_mem[8'h54] <= 8'h6a;
m11_mem[8'h55] <= 8'h61;
m11_mem[8'h56] <= 8'h7c;
m11_mem[8'h57] <= 8'h77;
m11_mem[8'h58] <= 8'h1e;
m11_mem[8'h59] <= 8'h15;
m11_mem[8'h5a] <= 8'h08;
m11_mem[8'h5b] <= 8'h03;
m11_mem[8'h5c] <= 8'h32;
m11_mem[8'h5d] <= 8'h39;
m11_mem[8'h5e] <= 8'h24;
m11_mem[8'h5f] <= 8'h2f;
m11_mem[8'h60] <= 8'h8d;
m11_mem[8'h61] <= 8'h86;
m11_mem[8'h62] <= 8'h9b;
m11_mem[8'h63] <= 8'h90;
m11_mem[8'h64] <= 8'ha1;
m11_mem[8'h65] <= 8'haa;
m11_mem[8'h66] <= 8'hb7;
m11_mem[8'h67] <= 8'hbc;
m11_mem[8'h68] <= 8'hd5;
m11_mem[8'h69] <= 8'hde;
m11_mem[8'h6a] <= 8'hc3;
m11_mem[8'h6b] <= 8'hc8;
m11_mem[8'h6c] <= 8'hf9;
m11_mem[8'h6d] <= 8'hf2;
m11_mem[8'h6e] <= 8'hef;
m11_mem[8'h6f] <= 8'he4;
m11_mem[8'h70] <= 8'h3d;
m11_mem[8'h71] <= 8'h36;
m11_mem[8'h72] <= 8'h2b;
m11_mem[8'h73] <= 8'h20;
m11_mem[8'h74] <= 8'h11;
m11_mem[8'h75] <= 8'h1a;
m11_mem[8'h76] <= 8'h07;
m11_mem[8'h77] <= 8'h0c;
m11_mem[8'h78] <= 8'h65;
m11_mem[8'h79] <= 8'h6e;
m11_mem[8'h7a] <= 8'h73;
m11_mem[8'h7b] <= 8'h78;
m11_mem[8'h7c] <= 8'h49;
m11_mem[8'h7d] <= 8'h42;
m11_mem[8'h7e] <= 8'h5f;
m11_mem[8'h7f] <= 8'h54;
m11_mem[8'h80] <= 8'hf7;
m11_mem[8'h81] <= 8'hfc;
m11_mem[8'h82] <= 8'he1;
m11_mem[8'h83] <= 8'hea;
m11_mem[8'h84] <= 8'hdb;
m11_mem[8'h85] <= 8'hd0;
m11_mem[8'h86] <= 8'hcd;
m11_mem[8'h87] <= 8'hc6;
m11_mem[8'h88] <= 8'haf;
m11_mem[8'h89] <= 8'ha4;
m11_mem[8'h8a] <= 8'hb9;
m11_mem[8'h8b] <= 8'hb2;
m11_mem[8'h8c] <= 8'h83;
m11_mem[8'h8d] <= 8'h88;
m11_mem[8'h8e] <= 8'h95;
m11_mem[8'h8f] <= 8'h9e;
m11_mem[8'h90] <= 8'h47;
m11_mem[8'h91] <= 8'h4c;
m11_mem[8'h92] <= 8'h51;
m11_mem[8'h93] <= 8'h5a;
m11_mem[8'h94] <= 8'h6b;
m11_mem[8'h95] <= 8'h60;
m11_mem[8'h96] <= 8'h7d;
m11_mem[8'h97] <= 8'h76;
m11_mem[8'h98] <= 8'h1f;
m11_mem[8'h99] <= 8'h14;
m11_mem[8'h9a] <= 8'h09;
m11_mem[8'h9b] <= 8'h02;
m11_mem[8'h9c] <= 8'h33;
m11_mem[8'h9d] <= 8'h38;
m11_mem[8'h9e] <= 8'h25;
m11_mem[8'h9f] <= 8'h2e;
m11_mem[8'ha0] <= 8'h8c;
m11_mem[8'ha1] <= 8'h87;
m11_mem[8'ha2] <= 8'h9a;
m11_mem[8'ha3] <= 8'h91;
m11_mem[8'ha4] <= 8'ha0;
m11_mem[8'ha5] <= 8'hab;
m11_mem[8'ha6] <= 8'hb6;
m11_mem[8'ha7] <= 8'hbd;
m11_mem[8'ha8] <= 8'hd4;
m11_mem[8'ha9] <= 8'hdf;
m11_mem[8'haa] <= 8'hc2;
m11_mem[8'hab] <= 8'hc9;
m11_mem[8'hac] <= 8'hf8;
m11_mem[8'had] <= 8'hf3;
m11_mem[8'hae] <= 8'hee;
m11_mem[8'haf] <= 8'he5;
m11_mem[8'hb0] <= 8'h3c;
m11_mem[8'hb1] <= 8'h37;
m11_mem[8'hb2] <= 8'h2a;
m11_mem[8'hb3] <= 8'h21;
m11_mem[8'hb4] <= 8'h10;
m11_mem[8'hb5] <= 8'h1b;
m11_mem[8'hb6] <= 8'h06;
m11_mem[8'hb7] <= 8'h0d;
m11_mem[8'hb8] <= 8'h64;
m11_mem[8'hb9] <= 8'h6f;
m11_mem[8'hba] <= 8'h72;
m11_mem[8'hbb] <= 8'h79;
m11_mem[8'hbc] <= 8'h48;
m11_mem[8'hbd] <= 8'h43;
m11_mem[8'hbe] <= 8'h5e;
m11_mem[8'hbf] <= 8'h55;
m11_mem[8'hc0] <= 8'h01;
m11_mem[8'hc1] <= 8'h0a;
m11_mem[8'hc2] <= 8'h17;
m11_mem[8'hc3] <= 8'h1c;
m11_mem[8'hc4] <= 8'h2d;
m11_mem[8'hc5] <= 8'h26;
m11_mem[8'hc6] <= 8'h3b;
m11_mem[8'hc7] <= 8'h30;
m11_mem[8'hc8] <= 8'h59;
m11_mem[8'hc9] <= 8'h52;
m11_mem[8'hca] <= 8'h4f;
m11_mem[8'hcb] <= 8'h44;
m11_mem[8'hcc] <= 8'h75;
m11_mem[8'hcd] <= 8'h7e;
m11_mem[8'hce] <= 8'h63;
m11_mem[8'hcf] <= 8'h68;
m11_mem[8'hd0] <= 8'hb1;
m11_mem[8'hd1] <= 8'hba;
m11_mem[8'hd2] <= 8'ha7;
m11_mem[8'hd3] <= 8'hac;
m11_mem[8'hd4] <= 8'h9d;
m11_mem[8'hd5] <= 8'h96;
m11_mem[8'hd6] <= 8'h8b;
m11_mem[8'hd7] <= 8'h80;
m11_mem[8'hd8] <= 8'he9;
m11_mem[8'hd9] <= 8'he2;
m11_mem[8'hda] <= 8'hff;
m11_mem[8'hdb] <= 8'hf4;
m11_mem[8'hdc] <= 8'hc5;
m11_mem[8'hdd] <= 8'hce;
m11_mem[8'hde] <= 8'hd3;
m11_mem[8'hdf] <= 8'hd8;
m11_mem[8'he0] <= 8'h7a;
m11_mem[8'he1] <= 8'h71;
m11_mem[8'he2] <= 8'h6c;
m11_mem[8'he3] <= 8'h67;
m11_mem[8'he4] <= 8'h56;
m11_mem[8'he5] <= 8'h5d;
m11_mem[8'he6] <= 8'h40;
m11_mem[8'he7] <= 8'h4b;
m11_mem[8'he8] <= 8'h22;
m11_mem[8'he9] <= 8'h29;
m11_mem[8'hea] <= 8'h34;
m11_mem[8'heb] <= 8'h3f;
m11_mem[8'hec] <= 8'h0e;
m11_mem[8'hed] <= 8'h05;
m11_mem[8'hee] <= 8'h18;
m11_mem[8'hef] <= 8'h13;
m11_mem[8'hf0] <= 8'hca;
m11_mem[8'hf1] <= 8'hc1;
m11_mem[8'hf2] <= 8'hdc;
m11_mem[8'hf3] <= 8'hd7;
m11_mem[8'hf4] <= 8'he6;
m11_mem[8'hf5] <= 8'hed;
m11_mem[8'hf6] <= 8'hf0;
m11_mem[8'hf7] <= 8'hfb;
m11_mem[8'hf8] <= 8'h92;
m11_mem[8'hf9] <= 8'h99;
m11_mem[8'hfa] <= 8'h84;
m11_mem[8'hfb] <= 8'h8f;
m11_mem[8'hfc] <= 8'hbe;
m11_mem[8'hfd] <= 8'hb5;
m11_mem[8'hfe] <= 8'ha8;
m11_mem[8'hff] <= 8'ha3;
end

endmodule
