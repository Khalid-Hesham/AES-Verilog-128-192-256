module M2 (
  input [7:0] in,
  output reg [7:0] out
);

reg [7:0] m2_mem [0:255] ;

always @(*) out = m2_mem[in];


initial begin
m2_mem[8'h00] <= 8'h00;
m2_mem[8'h01] <= 8'h02;
m2_mem[8'h02] <= 8'h04;
m2_mem[8'h03] <= 8'h06;
m2_mem[8'h04] <= 8'h08;
m2_mem[8'h05] <= 8'h0a;
m2_mem[8'h06] <= 8'h0c;
m2_mem[8'h07] <= 8'h0e;
m2_mem[8'h08] <= 8'h10;
m2_mem[8'h09] <= 8'h12;
m2_mem[8'h0a] <= 8'h14;
m2_mem[8'h0b] <= 8'h16;
m2_mem[8'h0c] <= 8'h18;
m2_mem[8'h0d] <= 8'h1a;
m2_mem[8'h0e] <= 8'h1c;
m2_mem[8'h0f] <= 8'h1e;
m2_mem[8'h10] <= 8'h20;
m2_mem[8'h11] <= 8'h22;
m2_mem[8'h12] <= 8'h24;
m2_mem[8'h13] <= 8'h26;
m2_mem[8'h14] <= 8'h28;
m2_mem[8'h15] <= 8'h2a;
m2_mem[8'h16] <= 8'h2c;
m2_mem[8'h17] <= 8'h2e;
m2_mem[8'h18] <= 8'h30;
m2_mem[8'h19] <= 8'h32;
m2_mem[8'h1a] <= 8'h34;
m2_mem[8'h1b] <= 8'h36;
m2_mem[8'h1c] <= 8'h38;
m2_mem[8'h1d] <= 8'h3a;
m2_mem[8'h1e] <= 8'h3c;
m2_mem[8'h1f] <= 8'h3e;
m2_mem[8'h20] <= 8'h40;
m2_mem[8'h21] <= 8'h42;
m2_mem[8'h22] <= 8'h44;
m2_mem[8'h23] <= 8'h46;
m2_mem[8'h24] <= 8'h48;
m2_mem[8'h25] <= 8'h4a;
m2_mem[8'h26] <= 8'h4c;
m2_mem[8'h27] <= 8'h4e;
m2_mem[8'h28] <= 8'h50;
m2_mem[8'h29] <= 8'h52;
m2_mem[8'h2a] <= 8'h54;
m2_mem[8'h2b] <= 8'h56;
m2_mem[8'h2c] <= 8'h58;
m2_mem[8'h2d] <= 8'h5a;
m2_mem[8'h2e] <= 8'h5c;
m2_mem[8'h2f] <= 8'h5e;
m2_mem[8'h30] <= 8'h60;
m2_mem[8'h31] <= 8'h62;
m2_mem[8'h32] <= 8'h64;
m2_mem[8'h33] <= 8'h66;
m2_mem[8'h34] <= 8'h68;
m2_mem[8'h35] <= 8'h6a;
m2_mem[8'h36] <= 8'h6c;
m2_mem[8'h37] <= 8'h6e;
m2_mem[8'h38] <= 8'h70;
m2_mem[8'h39] <= 8'h72;
m2_mem[8'h3a] <= 8'h74;
m2_mem[8'h3b] <= 8'h76;
m2_mem[8'h3c] <= 8'h78;
m2_mem[8'h3d] <= 8'h7a;
m2_mem[8'h3e] <= 8'h7c;
m2_mem[8'h3f] <= 8'h7e;
m2_mem[8'h40] <= 8'h80;
m2_mem[8'h41] <= 8'h82;
m2_mem[8'h42] <= 8'h84;
m2_mem[8'h43] <= 8'h86;
m2_mem[8'h44] <= 8'h88;
m2_mem[8'h45] <= 8'h8a;
m2_mem[8'h46] <= 8'h8c;
m2_mem[8'h47] <= 8'h8e;
m2_mem[8'h48] <= 8'h90;
m2_mem[8'h49] <= 8'h92;
m2_mem[8'h4a] <= 8'h94;
m2_mem[8'h4b] <= 8'h96;
m2_mem[8'h4c] <= 8'h98;
m2_mem[8'h4d] <= 8'h9a;
m2_mem[8'h4e] <= 8'h9c;
m2_mem[8'h4f] <= 8'h9e;
m2_mem[8'h50] <= 8'ha0;
m2_mem[8'h51] <= 8'ha2;
m2_mem[8'h52] <= 8'ha4;
m2_mem[8'h53] <= 8'ha6;
m2_mem[8'h54] <= 8'ha8;
m2_mem[8'h55] <= 8'haa;
m2_mem[8'h56] <= 8'hac;
m2_mem[8'h57] <= 8'hae;
m2_mem[8'h58] <= 8'hb0;
m2_mem[8'h59] <= 8'hb2;
m2_mem[8'h5a] <= 8'hb4;
m2_mem[8'h5b] <= 8'hb6;
m2_mem[8'h5c] <= 8'hb8;
m2_mem[8'h5d] <= 8'hba;
m2_mem[8'h5e] <= 8'hbc;
m2_mem[8'h5f] <= 8'hbe;
m2_mem[8'h60] <= 8'hc0;
m2_mem[8'h61] <= 8'hc2;
m2_mem[8'h62] <= 8'hc4;
m2_mem[8'h63] <= 8'hc6;
m2_mem[8'h64] <= 8'hc8;
m2_mem[8'h65] <= 8'hca;
m2_mem[8'h66] <= 8'hcc;
m2_mem[8'h67] <= 8'hce;
m2_mem[8'h68] <= 8'hd0;
m2_mem[8'h69] <= 8'hd2;
m2_mem[8'h6a] <= 8'hd4;
m2_mem[8'h6b] <= 8'hd6;
m2_mem[8'h6c] <= 8'hd8;
m2_mem[8'h6d] <= 8'hda;
m2_mem[8'h6e] <= 8'hdc;
m2_mem[8'h6f] <= 8'hde;
m2_mem[8'h70] <= 8'he0;
m2_mem[8'h71] <= 8'he2;
m2_mem[8'h72] <= 8'he4;
m2_mem[8'h73] <= 8'he6;
m2_mem[8'h74] <= 8'he8;
m2_mem[8'h75] <= 8'hea;
m2_mem[8'h76] <= 8'hec;
m2_mem[8'h77] <= 8'hee;
m2_mem[8'h78] <= 8'hf0;
m2_mem[8'h79] <= 8'hf2;
m2_mem[8'h7a] <= 8'hf4;
m2_mem[8'h7b] <= 8'hf6;
m2_mem[8'h7c] <= 8'hf8;
m2_mem[8'h7d] <= 8'hfa;
m2_mem[8'h7e] <= 8'hfc;
m2_mem[8'h7f] <= 8'hfe;
m2_mem[8'h80] <= 8'h1b;
m2_mem[8'h81] <= 8'h19;
m2_mem[8'h82] <= 8'h1f;
m2_mem[8'h83] <= 8'h1d;
m2_mem[8'h84] <= 8'h13;
m2_mem[8'h85] <= 8'h11;
m2_mem[8'h86] <= 8'h17;
m2_mem[8'h87] <= 8'h15;
m2_mem[8'h88] <= 8'h0b;
m2_mem[8'h89] <= 8'h09;
m2_mem[8'h8a] <= 8'h0f;
m2_mem[8'h8b] <= 8'h0d;
m2_mem[8'h8c] <= 8'h03;
m2_mem[8'h8d] <= 8'h01;
m2_mem[8'h8e] <= 8'h07;
m2_mem[8'h8f] <= 8'h05;
m2_mem[8'h90] <= 8'h3b;
m2_mem[8'h91] <= 8'h39;
m2_mem[8'h92] <= 8'h3f;
m2_mem[8'h93] <= 8'h3d;
m2_mem[8'h94] <= 8'h33;
m2_mem[8'h95] <= 8'h31;
m2_mem[8'h96] <= 8'h37;
m2_mem[8'h97] <= 8'h35;
m2_mem[8'h98] <= 8'h2b;
m2_mem[8'h99] <= 8'h29;
m2_mem[8'h9a] <= 8'h2f;
m2_mem[8'h9b] <= 8'h2d;
m2_mem[8'h9c] <= 8'h23;
m2_mem[8'h9d] <= 8'h21;
m2_mem[8'h9e] <= 8'h27;
m2_mem[8'h9f] <= 8'h25;
m2_mem[8'ha0] <= 8'h5b;
m2_mem[8'ha1] <= 8'h59;
m2_mem[8'ha2] <= 8'h5f;
m2_mem[8'ha3] <= 8'h5d;
m2_mem[8'ha4] <= 8'h53;
m2_mem[8'ha5] <= 8'h51;
m2_mem[8'ha6] <= 8'h57;
m2_mem[8'ha7] <= 8'h55;
m2_mem[8'ha8] <= 8'h4b;
m2_mem[8'ha9] <= 8'h49;
m2_mem[8'haa] <= 8'h4f;
m2_mem[8'hab] <= 8'h4d;
m2_mem[8'hac] <= 8'h43;
m2_mem[8'had] <= 8'h41;
m2_mem[8'hae] <= 8'h47;
m2_mem[8'haf] <= 8'h45;
m2_mem[8'hb0] <= 8'h7b;
m2_mem[8'hb1] <= 8'h79;
m2_mem[8'hb2] <= 8'h7f;
m2_mem[8'hb3] <= 8'h7d;
m2_mem[8'hb4] <= 8'h73;
m2_mem[8'hb5] <= 8'h71;
m2_mem[8'hb6] <= 8'h77;
m2_mem[8'hb7] <= 8'h75;
m2_mem[8'hb8] <= 8'h6b;
m2_mem[8'hb9] <= 8'h69;
m2_mem[8'hba] <= 8'h6f;
m2_mem[8'hbb] <= 8'h6d;
m2_mem[8'hbc] <= 8'h63;
m2_mem[8'hbd] <= 8'h61;
m2_mem[8'hbe] <= 8'h67;
m2_mem[8'hbf] <= 8'h65;
m2_mem[8'hc0] <= 8'h9b;
m2_mem[8'hc1] <= 8'h99;
m2_mem[8'hc2] <= 8'h9f;
m2_mem[8'hc3] <= 8'h9d;
m2_mem[8'hc4] <= 8'h93;
m2_mem[8'hc5] <= 8'h91;
m2_mem[8'hc6] <= 8'h97;
m2_mem[8'hc7] <= 8'h95;
m2_mem[8'hc8] <= 8'h8b;
m2_mem[8'hc9] <= 8'h89;
m2_mem[8'hca] <= 8'h8f;
m2_mem[8'hcb] <= 8'h8d;
m2_mem[8'hcc] <= 8'h83;
m2_mem[8'hcd] <= 8'h81;
m2_mem[8'hce] <= 8'h87;
m2_mem[8'hcf] <= 8'h85;
m2_mem[8'hd0] <= 8'hbb;
m2_mem[8'hd1] <= 8'hb9;
m2_mem[8'hd2] <= 8'hbf;
m2_mem[8'hd3] <= 8'hbd;
m2_mem[8'hd4] <= 8'hb3;
m2_mem[8'hd5] <= 8'hb1;
m2_mem[8'hd6] <= 8'hb7;
m2_mem[8'hd7] <= 8'hb5;
m2_mem[8'hd8] <= 8'hab;
m2_mem[8'hd9] <= 8'ha9;
m2_mem[8'hda] <= 8'haf;
m2_mem[8'hdb] <= 8'had;
m2_mem[8'hdc] <= 8'ha3;
m2_mem[8'hdd] <= 8'ha1;
m2_mem[8'hde] <= 8'ha7;
m2_mem[8'hdf] <= 8'ha5;
m2_mem[8'he0] <= 8'hdb;
m2_mem[8'he1] <= 8'hd9;
m2_mem[8'he2] <= 8'hdf;
m2_mem[8'he3] <= 8'hdd;
m2_mem[8'he4] <= 8'hd3;
m2_mem[8'he5] <= 8'hd1;
m2_mem[8'he6] <= 8'hd7;
m2_mem[8'he7] <= 8'hd5;
m2_mem[8'he8] <= 8'hcb;
m2_mem[8'he9] <= 8'hc9;
m2_mem[8'hea] <= 8'hcf;
m2_mem[8'heb] <= 8'hcd;
m2_mem[8'hec] <= 8'hc3;
m2_mem[8'hed] <= 8'hc1;
m2_mem[8'hee] <= 8'hc7;
m2_mem[8'hef] <= 8'hc5;
m2_mem[8'hf0] <= 8'hfb;
m2_mem[8'hf1] <= 8'hf9;
m2_mem[8'hf2] <= 8'hff;
m2_mem[8'hf3] <= 8'hfd;
m2_mem[8'hf4] <= 8'hf3;
m2_mem[8'hf5] <= 8'hf1;
m2_mem[8'hf6] <= 8'hf7;
m2_mem[8'hf7] <= 8'hf5;
m2_mem[8'hf8] <= 8'heb;
m2_mem[8'hf9] <= 8'he9;
m2_mem[8'hfa] <= 8'hef;
m2_mem[8'hfb] <= 8'hed;
m2_mem[8'hfc] <= 8'he3;
m2_mem[8'hfd] <= 8'he1;
m2_mem[8'hfe] <= 8'he7;
m2_mem[8'hff] <= 8'he5;  
end


endmodule
