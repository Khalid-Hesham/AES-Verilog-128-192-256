module inv_sbox (
  input [7:0] in,
  output reg [7:0] out
);

reg [7:0] isb_mem [0:255];

always @(*) out = isb_mem[in];

initial begin
isb_mem[8'h00] <= 8'h52;
isb_mem[8'h01] <= 8'h09;
isb_mem[8'h02] <= 8'h6a;
isb_mem[8'h03] <= 8'hd5;
isb_mem[8'h04] <= 8'h30;
isb_mem[8'h05] <= 8'h36;
isb_mem[8'h06] <= 8'ha5;
isb_mem[8'h07] <= 8'h38;
isb_mem[8'h08] <= 8'hbf;
isb_mem[8'h09] <= 8'h40;
isb_mem[8'h0a] <= 8'ha3;
isb_mem[8'h0b] <= 8'h9e;
isb_mem[8'h0c] <= 8'h81;
isb_mem[8'h0d] <= 8'hf3;
isb_mem[8'h0e] <= 8'hd7;
isb_mem[8'h0f] <= 8'hfb;
isb_mem[8'h10] <= 8'h7c;
isb_mem[8'h11] <= 8'he3;
isb_mem[8'h12] <= 8'h39;
isb_mem[8'h13] <= 8'h82;
isb_mem[8'h14] <= 8'h9b;
isb_mem[8'h15] <= 8'h2f;
isb_mem[8'h16] <= 8'hff;
isb_mem[8'h17] <= 8'h87;
isb_mem[8'h18] <= 8'h34;
isb_mem[8'h19] <= 8'h8e;
isb_mem[8'h1a] <= 8'h43;
isb_mem[8'h1b] <= 8'h44;
isb_mem[8'h1c] <= 8'hc4;
isb_mem[8'h1d] <= 8'hde;
isb_mem[8'h1e] <= 8'he9;
isb_mem[8'h1f] <= 8'hcb;
isb_mem[8'h20] <= 8'h54;
isb_mem[8'h21] <= 8'h7b;
isb_mem[8'h22] <= 8'h94;
isb_mem[8'h23] <= 8'h32;
isb_mem[8'h24] <= 8'ha6;
isb_mem[8'h25] <= 8'hc2;
isb_mem[8'h26] <= 8'h23;
isb_mem[8'h27] <= 8'h3d;
isb_mem[8'h28] <= 8'hee;
isb_mem[8'h29] <= 8'h4c;
isb_mem[8'h2a] <= 8'h95;
isb_mem[8'h2b] <= 8'h0b;
isb_mem[8'h2c] <= 8'h42;
isb_mem[8'h2d] <= 8'hfa;
isb_mem[8'h2e] <= 8'hc3;
isb_mem[8'h2f] <= 8'h4e;
isb_mem[8'h30] <= 8'h08;
isb_mem[8'h31] <= 8'h2e;
isb_mem[8'h32] <= 8'ha1;
isb_mem[8'h33] <= 8'h66;
isb_mem[8'h34] <= 8'h28;
isb_mem[8'h35] <= 8'hd9;
isb_mem[8'h36] <= 8'h24;
isb_mem[8'h37] <= 8'hb2;
isb_mem[8'h38] <= 8'h76;
isb_mem[8'h39] <= 8'h5b;
isb_mem[8'h3a] <= 8'ha2;
isb_mem[8'h3b] <= 8'h49;
isb_mem[8'h3c] <= 8'h6d;
isb_mem[8'h3d] <= 8'h8b;
isb_mem[8'h3e] <= 8'hd1;
isb_mem[8'h3f] <= 8'h25;
isb_mem[8'h40] <= 8'h72;
isb_mem[8'h41] <= 8'hf8;
isb_mem[8'h42] <= 8'hf6;
isb_mem[8'h43] <= 8'h64;
isb_mem[8'h44] <= 8'h86;
isb_mem[8'h45] <= 8'h68;
isb_mem[8'h46] <= 8'h98;
isb_mem[8'h47] <= 8'h16;
isb_mem[8'h48] <= 8'hd4;
isb_mem[8'h49] <= 8'ha4;
isb_mem[8'h4a] <= 8'h5c;
isb_mem[8'h4b] <= 8'hcc;
isb_mem[8'h4c] <= 8'h5d;
isb_mem[8'h4d] <= 8'h65;
isb_mem[8'h4e] <= 8'hb6;
isb_mem[8'h4f] <= 8'h92;
isb_mem[8'h50] <= 8'h6c;
isb_mem[8'h51] <= 8'h70;
isb_mem[8'h52] <= 8'h48;
isb_mem[8'h53] <= 8'h50;
isb_mem[8'h54] <= 8'hfd;
isb_mem[8'h55] <= 8'hed;
isb_mem[8'h56] <= 8'hb9;
isb_mem[8'h57] <= 8'hda;
isb_mem[8'h58] <= 8'h5e;
isb_mem[8'h59] <= 8'h15;
isb_mem[8'h5a] <= 8'h46;
isb_mem[8'h5b] <= 8'h57;
isb_mem[8'h5c] <= 8'ha7;
isb_mem[8'h5d] <= 8'h8d;
isb_mem[8'h5e] <= 8'h9d;
isb_mem[8'h5f] <= 8'h84;
isb_mem[8'h60] <= 8'h90;
isb_mem[8'h61] <= 8'hd8;
isb_mem[8'h62] <= 8'hab;
isb_mem[8'h63] <= 8'h00;
isb_mem[8'h64] <= 8'h8c;
isb_mem[8'h65] <= 8'hbc;
isb_mem[8'h66] <= 8'hd3;
isb_mem[8'h67] <= 8'h0a;
isb_mem[8'h68] <= 8'hf7;
isb_mem[8'h69] <= 8'he4;
isb_mem[8'h6a] <= 8'h58;
isb_mem[8'h6b] <= 8'h05;
isb_mem[8'h6c] <= 8'hb8;
isb_mem[8'h6d] <= 8'hb3;
isb_mem[8'h6e] <= 8'h45;
isb_mem[8'h6f] <= 8'h06;
isb_mem[8'h70] <= 8'hd0;
isb_mem[8'h71] <= 8'h2c;
isb_mem[8'h72] <= 8'h1e;
isb_mem[8'h73] <= 8'h8f;
isb_mem[8'h74] <= 8'hca;
isb_mem[8'h75] <= 8'h3f;
isb_mem[8'h76] <= 8'h0f;
isb_mem[8'h77] <= 8'h02;
isb_mem[8'h78] <= 8'hc1;
isb_mem[8'h79] <= 8'haf;
isb_mem[8'h7a] <= 8'hbd;
isb_mem[8'h7b] <= 8'h03;
isb_mem[8'h7c] <= 8'h01;
isb_mem[8'h7d] <= 8'h13;
isb_mem[8'h7e] <= 8'h8a;
isb_mem[8'h7f] <= 8'h6b;
isb_mem[8'h80] <= 8'h3a;
isb_mem[8'h81] <= 8'h91;
isb_mem[8'h82] <= 8'h11;
isb_mem[8'h83] <= 8'h41;
isb_mem[8'h84] <= 8'h4f;
isb_mem[8'h85] <= 8'h67;
isb_mem[8'h86] <= 8'hdc;
isb_mem[8'h87] <= 8'hea;
isb_mem[8'h88] <= 8'h97;
isb_mem[8'h89] <= 8'hf2;
isb_mem[8'h8a] <= 8'hcf;
isb_mem[8'h8b] <= 8'hce;
isb_mem[8'h8c] <= 8'hf0;
isb_mem[8'h8d] <= 8'hb4;
isb_mem[8'h8e] <= 8'he6;
isb_mem[8'h8f] <= 8'h73;
isb_mem[8'h90] <= 8'h96;
isb_mem[8'h91] <= 8'hac;
isb_mem[8'h92] <= 8'h74;
isb_mem[8'h93] <= 8'h22;
isb_mem[8'h94] <= 8'he7;
isb_mem[8'h95] <= 8'had;
isb_mem[8'h96] <= 8'h35;
isb_mem[8'h97] <= 8'h85;
isb_mem[8'h98] <= 8'he2;
isb_mem[8'h99] <= 8'hf9;
isb_mem[8'h9a] <= 8'h37;
isb_mem[8'h9b] <= 8'he8;
isb_mem[8'h9c] <= 8'h1c;
isb_mem[8'h9d] <= 8'h75;
isb_mem[8'h9e] <= 8'hdf;
isb_mem[8'h9f] <= 8'h6e;
isb_mem[8'ha0] <= 8'h47;
isb_mem[8'ha1] <= 8'hf1;
isb_mem[8'ha2] <= 8'h1a;
isb_mem[8'ha3] <= 8'h71;
isb_mem[8'ha4] <= 8'h1d;
isb_mem[8'ha5] <= 8'h29;
isb_mem[8'ha6] <= 8'hc5;
isb_mem[8'ha7] <= 8'h89;
isb_mem[8'ha8] <= 8'h6f;
isb_mem[8'ha9] <= 8'hb7;
isb_mem[8'haa] <= 8'h62;
isb_mem[8'hab] <= 8'h0e;
isb_mem[8'hac] <= 8'haa;
isb_mem[8'had] <= 8'h18;
isb_mem[8'hae] <= 8'hbe;
isb_mem[8'haf] <= 8'h1b;
isb_mem[8'hb0] <= 8'hfc;
isb_mem[8'hb1] <= 8'h56;
isb_mem[8'hb2] <= 8'h3e;
isb_mem[8'hb3] <= 8'h4b;
isb_mem[8'hb4] <= 8'hc6;
isb_mem[8'hb5] <= 8'hd2;
isb_mem[8'hb6] <= 8'h79;
isb_mem[8'hb7] <= 8'h20;
isb_mem[8'hb8] <= 8'h9a;
isb_mem[8'hb9] <= 8'hdb;
isb_mem[8'hba] <= 8'hc0;
isb_mem[8'hbb] <= 8'hfe;
isb_mem[8'hbc] <= 8'h78;
isb_mem[8'hbd] <= 8'hcd;
isb_mem[8'hbe] <= 8'h5a;
isb_mem[8'hbf] <= 8'hf4;
isb_mem[8'hc0] <= 8'h1f;
isb_mem[8'hc1] <= 8'hdd;
isb_mem[8'hc2] <= 8'ha8;
isb_mem[8'hc3] <= 8'h33;
isb_mem[8'hc4] <= 8'h88;
isb_mem[8'hc5] <= 8'h07;
isb_mem[8'hc6] <= 8'hc7;
isb_mem[8'hc7] <= 8'h31;
isb_mem[8'hc8] <= 8'hb1;
isb_mem[8'hc9] <= 8'h12;
isb_mem[8'hca] <= 8'h10;
isb_mem[8'hcb] <= 8'h59;
isb_mem[8'hcc] <= 8'h27;
isb_mem[8'hcd] <= 8'h80;
isb_mem[8'hce] <= 8'hec;
isb_mem[8'hcf] <= 8'h5f;
isb_mem[8'hd0] <= 8'h60;
isb_mem[8'hd1] <= 8'h51;
isb_mem[8'hd2] <= 8'h7f;
isb_mem[8'hd3] <= 8'ha9;
isb_mem[8'hd4] <= 8'h19;
isb_mem[8'hd5] <= 8'hb5;
isb_mem[8'hd6] <= 8'h4a;
isb_mem[8'hd7] <= 8'h0d;
isb_mem[8'hd8] <= 8'h2d;
isb_mem[8'hd9] <= 8'he5;
isb_mem[8'hda] <= 8'h7a;
isb_mem[8'hdb] <= 8'h9f;
isb_mem[8'hdc] <= 8'h93;
isb_mem[8'hdd] <= 8'hc9;
isb_mem[8'hde] <= 8'h9c;
isb_mem[8'hdf] <= 8'hef;
isb_mem[8'he0] <= 8'ha0;
isb_mem[8'he1] <= 8'he0;
isb_mem[8'he2] <= 8'h3b;
isb_mem[8'he3] <= 8'h4d;
isb_mem[8'he4] <= 8'hae;
isb_mem[8'he5] <= 8'h2a;
isb_mem[8'he6] <= 8'hf5;
isb_mem[8'he7] <= 8'hb0;
isb_mem[8'he8] <= 8'hc8;
isb_mem[8'he9] <= 8'heb;
isb_mem[8'hea] <= 8'hbb;
isb_mem[8'heb] <= 8'h3c;
isb_mem[8'hec] <= 8'h83;
isb_mem[8'hed] <= 8'h53;
isb_mem[8'hee] <= 8'h99;
isb_mem[8'hef] <= 8'h61;
isb_mem[8'hf0] <= 8'h17;
isb_mem[8'hf1] <= 8'h2b;
isb_mem[8'hf2] <= 8'h04;
isb_mem[8'hf3] <= 8'h7e;
isb_mem[8'hf4] <= 8'hba;
isb_mem[8'hf5] <= 8'h77;
isb_mem[8'hf6] <= 8'hd6;
isb_mem[8'hf7] <= 8'h26;
isb_mem[8'hf8] <= 8'he1;
isb_mem[8'hf9] <= 8'h69;
isb_mem[8'hfa] <= 8'h14;
isb_mem[8'hfb] <= 8'h63;
isb_mem[8'hfc] <= 8'h55;
isb_mem[8'hfd] <= 8'h21;
isb_mem[8'hfe] <= 8'h0c;
isb_mem[8'hff] <= 8'h7d;
end



endmodule 
