module M9 (
  input [7:0] in,
  output reg [7:0] out
);

reg [7:0] m9_mem [0:255]; 

always @(*) out = m9_mem[in];

initial begin
m9_mem[8'h00] <= 8'h00;
m9_mem[8'h01] <= 8'h09;
m9_mem[8'h02] <= 8'h12;
m9_mem[8'h03] <= 8'h1b;
m9_mem[8'h04] <= 8'h24;
m9_mem[8'h05] <= 8'h2d;
m9_mem[8'h06] <= 8'h36;
m9_mem[8'h07] <= 8'h3f;
m9_mem[8'h08] <= 8'h48;
m9_mem[8'h09] <= 8'h41;
m9_mem[8'h0a] <= 8'h5a;
m9_mem[8'h0b] <= 8'h53;
m9_mem[8'h0c] <= 8'h6c;
m9_mem[8'h0d] <= 8'h65;
m9_mem[8'h0e] <= 8'h7e;
m9_mem[8'h0f] <= 8'h77;
m9_mem[8'h10] <= 8'h90;
m9_mem[8'h11] <= 8'h99;
m9_mem[8'h12] <= 8'h82;
m9_mem[8'h13] <= 8'h8b;
m9_mem[8'h14] <= 8'hb4;
m9_mem[8'h15] <= 8'hbd;
m9_mem[8'h16] <= 8'ha6;
m9_mem[8'h17] <= 8'haf;
m9_mem[8'h18] <= 8'hd8;
m9_mem[8'h19] <= 8'hd1;
m9_mem[8'h1a] <= 8'hca;
m9_mem[8'h1b] <= 8'hc3;
m9_mem[8'h1c] <= 8'hfc;
m9_mem[8'h1d] <= 8'hf5;
m9_mem[8'h1e] <= 8'hee;
m9_mem[8'h1f] <= 8'he7;
m9_mem[8'h20] <= 8'h3b;
m9_mem[8'h21] <= 8'h32;
m9_mem[8'h22] <= 8'h29;
m9_mem[8'h23] <= 8'h20;
m9_mem[8'h24] <= 8'h1f;
m9_mem[8'h25] <= 8'h16;
m9_mem[8'h26] <= 8'h0d;
m9_mem[8'h27] <= 8'h04;
m9_mem[8'h28] <= 8'h73;
m9_mem[8'h29] <= 8'h7a;
m9_mem[8'h2a] <= 8'h61;
m9_mem[8'h2b] <= 8'h68;
m9_mem[8'h2c] <= 8'h57;
m9_mem[8'h2d] <= 8'h5e;
m9_mem[8'h2e] <= 8'h45;
m9_mem[8'h2f] <= 8'h4c;
m9_mem[8'h30] <= 8'hab;
m9_mem[8'h31] <= 8'ha2;
m9_mem[8'h32] <= 8'hb9;
m9_mem[8'h33] <= 8'hb0;
m9_mem[8'h34] <= 8'h8f;
m9_mem[8'h35] <= 8'h86;
m9_mem[8'h36] <= 8'h9d;
m9_mem[8'h37] <= 8'h94;
m9_mem[8'h38] <= 8'he3;
m9_mem[8'h39] <= 8'hea;
m9_mem[8'h3a] <= 8'hf1;
m9_mem[8'h3b] <= 8'hf8;
m9_mem[8'h3c] <= 8'hc7;
m9_mem[8'h3d] <= 8'hce;
m9_mem[8'h3e] <= 8'hd5;
m9_mem[8'h3f] <= 8'hdc;
m9_mem[8'h40] <= 8'h76;
m9_mem[8'h41] <= 8'h7f;
m9_mem[8'h42] <= 8'h64;
m9_mem[8'h43] <= 8'h6d;
m9_mem[8'h44] <= 8'h52;
m9_mem[8'h45] <= 8'h5b;
m9_mem[8'h46] <= 8'h40;
m9_mem[8'h47] <= 8'h49;
m9_mem[8'h48] <= 8'h3e;
m9_mem[8'h49] <= 8'h37;
m9_mem[8'h4a] <= 8'h2c;
m9_mem[8'h4b] <= 8'h25;
m9_mem[8'h4c] <= 8'h1a;
m9_mem[8'h4d] <= 8'h13;
m9_mem[8'h4e] <= 8'h08;
m9_mem[8'h4f] <= 8'h01;
m9_mem[8'h50] <= 8'he6;
m9_mem[8'h51] <= 8'hef;
m9_mem[8'h52] <= 8'hf4;
m9_mem[8'h53] <= 8'hfd;
m9_mem[8'h54] <= 8'hc2;
m9_mem[8'h55] <= 8'hcb;
m9_mem[8'h56] <= 8'hd0;
m9_mem[8'h57] <= 8'hd9;
m9_mem[8'h58] <= 8'hae;
m9_mem[8'h59] <= 8'ha7;
m9_mem[8'h5a] <= 8'hbc;
m9_mem[8'h5b] <= 8'hb5;
m9_mem[8'h5c] <= 8'h8a;
m9_mem[8'h5d] <= 8'h83;
m9_mem[8'h5e] <= 8'h98;
m9_mem[8'h5f] <= 8'h91;
m9_mem[8'h60] <= 8'h4d;
m9_mem[8'h61] <= 8'h44;
m9_mem[8'h62] <= 8'h5f;
m9_mem[8'h63] <= 8'h56;
m9_mem[8'h64] <= 8'h69;
m9_mem[8'h65] <= 8'h60;
m9_mem[8'h66] <= 8'h7b;
m9_mem[8'h67] <= 8'h72;
m9_mem[8'h68] <= 8'h05;
m9_mem[8'h69] <= 8'h0c;
m9_mem[8'h6a] <= 8'h17;
m9_mem[8'h6b] <= 8'h1e;
m9_mem[8'h6c] <= 8'h21;
m9_mem[8'h6d] <= 8'h28;
m9_mem[8'h6e] <= 8'h33;
m9_mem[8'h6f] <= 8'h3a;
m9_mem[8'h70] <= 8'hdd;
m9_mem[8'h71] <= 8'hd4;
m9_mem[8'h72] <= 8'hcf;
m9_mem[8'h73] <= 8'hc6;
m9_mem[8'h74] <= 8'hf9;
m9_mem[8'h75] <= 8'hf0;
m9_mem[8'h76] <= 8'heb;
m9_mem[8'h77] <= 8'he2;
m9_mem[8'h78] <= 8'h95;
m9_mem[8'h79] <= 8'h9c;
m9_mem[8'h7a] <= 8'h87;
m9_mem[8'h7b] <= 8'h8e;
m9_mem[8'h7c] <= 8'hb1;
m9_mem[8'h7d] <= 8'hb8;
m9_mem[8'h7e] <= 8'ha3;
m9_mem[8'h7f] <= 8'haa;
m9_mem[8'h80] <= 8'hec;
m9_mem[8'h81] <= 8'he5;
m9_mem[8'h82] <= 8'hfe;
m9_mem[8'h83] <= 8'hf7;
m9_mem[8'h84] <= 8'hc8;
m9_mem[8'h85] <= 8'hc1;
m9_mem[8'h86] <= 8'hda;
m9_mem[8'h87] <= 8'hd3;
m9_mem[8'h88] <= 8'ha4;
m9_mem[8'h89] <= 8'had;
m9_mem[8'h8a] <= 8'hb6;
m9_mem[8'h8b] <= 8'hbf;
m9_mem[8'h8c] <= 8'h80;
m9_mem[8'h8d] <= 8'h89;
m9_mem[8'h8e] <= 8'h92;
m9_mem[8'h8f] <= 8'h9b;
m9_mem[8'h90] <= 8'h7c;
m9_mem[8'h91] <= 8'h75;
m9_mem[8'h92] <= 8'h6e;
m9_mem[8'h93] <= 8'h67;
m9_mem[8'h94] <= 8'h58;
m9_mem[8'h95] <= 8'h51;
m9_mem[8'h96] <= 8'h4a;
m9_mem[8'h97] <= 8'h43;
m9_mem[8'h98] <= 8'h34;
m9_mem[8'h99] <= 8'h3d;
m9_mem[8'h9a] <= 8'h26;
m9_mem[8'h9b] <= 8'h2f;
m9_mem[8'h9c] <= 8'h10;
m9_mem[8'h9d] <= 8'h19;
m9_mem[8'h9e] <= 8'h02;
m9_mem[8'h9f] <= 8'h0b;
m9_mem[8'ha0] <= 8'hd7;
m9_mem[8'ha1] <= 8'hde;
m9_mem[8'ha2] <= 8'hc5;
m9_mem[8'ha3] <= 8'hcc;
m9_mem[8'ha4] <= 8'hf3;
m9_mem[8'ha5] <= 8'hfa;
m9_mem[8'ha6] <= 8'he1;
m9_mem[8'ha7] <= 8'he8;
m9_mem[8'ha8] <= 8'h9f;
m9_mem[8'ha9] <= 8'h96;
m9_mem[8'haa] <= 8'h8d;
m9_mem[8'hab] <= 8'h84;
m9_mem[8'hac] <= 8'hbb;
m9_mem[8'had] <= 8'hb2;
m9_mem[8'hae] <= 8'ha9;
m9_mem[8'haf] <= 8'ha0;
m9_mem[8'hb0] <= 8'h47;
m9_mem[8'hb1] <= 8'h4e;
m9_mem[8'hb2] <= 8'h55;
m9_mem[8'hb3] <= 8'h5c;
m9_mem[8'hb4] <= 8'h63;
m9_mem[8'hb5] <= 8'h6a;
m9_mem[8'hb6] <= 8'h71;
m9_mem[8'hb7] <= 8'h78;
m9_mem[8'hb8] <= 8'h0f;
m9_mem[8'hb9] <= 8'h06;
m9_mem[8'hba] <= 8'h1d;
m9_mem[8'hbb] <= 8'h14;
m9_mem[8'hbc] <= 8'h2b;
m9_mem[8'hbd] <= 8'h22;
m9_mem[8'hbe] <= 8'h39;
m9_mem[8'hbf] <= 8'h30;
m9_mem[8'hc0] <= 8'h9a;
m9_mem[8'hc1] <= 8'h93;
m9_mem[8'hc2] <= 8'h88;
m9_mem[8'hc3] <= 8'h81;
m9_mem[8'hc4] <= 8'hbe;
m9_mem[8'hc5] <= 8'hb7;
m9_mem[8'hc6] <= 8'hac;
m9_mem[8'hc7] <= 8'ha5;
m9_mem[8'hc8] <= 8'hd2;
m9_mem[8'hc9] <= 8'hdb;
m9_mem[8'hca] <= 8'hc0;
m9_mem[8'hcb] <= 8'hc9;
m9_mem[8'hcc] <= 8'hf6;
m9_mem[8'hcd] <= 8'hff;
m9_mem[8'hce] <= 8'he4;
m9_mem[8'hcf] <= 8'hed;
m9_mem[8'hd0] <= 8'h0a;
m9_mem[8'hd1] <= 8'h03;
m9_mem[8'hd2] <= 8'h18;
m9_mem[8'hd3] <= 8'h11;
m9_mem[8'hd4] <= 8'h2e;
m9_mem[8'hd5] <= 8'h27;
m9_mem[8'hd6] <= 8'h3c;
m9_mem[8'hd7] <= 8'h35;
m9_mem[8'hd8] <= 8'h42;
m9_mem[8'hd9] <= 8'h4b;
m9_mem[8'hda] <= 8'h50;
m9_mem[8'hdb] <= 8'h59;
m9_mem[8'hdc] <= 8'h66;
m9_mem[8'hdd] <= 8'h6f;
m9_mem[8'hde] <= 8'h74;
m9_mem[8'hdf] <= 8'h7d;
m9_mem[8'he0] <= 8'ha1;
m9_mem[8'he1] <= 8'ha8;
m9_mem[8'he2] <= 8'hb3;
m9_mem[8'he3] <= 8'hba;
m9_mem[8'he4] <= 8'h85;
m9_mem[8'he5] <= 8'h8c;
m9_mem[8'he6] <= 8'h97;
m9_mem[8'he7] <= 8'h9e;
m9_mem[8'he8] <= 8'he9;
m9_mem[8'he9] <= 8'he0;
m9_mem[8'hea] <= 8'hfb;
m9_mem[8'heb] <= 8'hf2;
m9_mem[8'hec] <= 8'hcd;
m9_mem[8'hed] <= 8'hc4;
m9_mem[8'hee] <= 8'hdf;
m9_mem[8'hef] <= 8'hd6;
m9_mem[8'hf0] <= 8'h31;
m9_mem[8'hf1] <= 8'h38;
m9_mem[8'hf2] <= 8'h23;
m9_mem[8'hf3] <= 8'h2a;
m9_mem[8'hf4] <= 8'h15;
m9_mem[8'hf5] <= 8'h1c;
m9_mem[8'hf6] <= 8'h07;
m9_mem[8'hf7] <= 8'h0e;
m9_mem[8'hf8] <= 8'h79;
m9_mem[8'hf9] <= 8'h70;
m9_mem[8'hfa] <= 8'h6b;
m9_mem[8'hfb] <= 8'h62;
m9_mem[8'hfc] <= 8'h5d;
m9_mem[8'hfd] <= 8'h54;
m9_mem[8'hfe] <= 8'h4f;
m9_mem[8'hff] <= 8'h46;
end


endmodule
