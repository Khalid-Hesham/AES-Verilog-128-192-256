module M14 (
  input [7:0] in,
  output reg [7:0] out
);

reg [7:0] m14_mem [0:255];

always @(*) out = m14_mem[in];

initial begin
m14_mem[8'h00] <= 8'h00;
m14_mem[8'h01] <= 8'h0e;
m14_mem[8'h02] <= 8'h1c;
m14_mem[8'h03] <= 8'h12;
m14_mem[8'h04] <= 8'h38;
m14_mem[8'h05] <= 8'h36;
m14_mem[8'h06] <= 8'h24;
m14_mem[8'h07] <= 8'h2a;
m14_mem[8'h08] <= 8'h70;
m14_mem[8'h09] <= 8'h7e;
m14_mem[8'h0a] <= 8'h6c;
m14_mem[8'h0b] <= 8'h62;
m14_mem[8'h0c] <= 8'h48;
m14_mem[8'h0d] <= 8'h46;
m14_mem[8'h0e] <= 8'h54;
m14_mem[8'h0f] <= 8'h5a;
m14_mem[8'h10] <= 8'he0;
m14_mem[8'h11] <= 8'hee;
m14_mem[8'h12] <= 8'hfc;
m14_mem[8'h13] <= 8'hf2;
m14_mem[8'h14] <= 8'hd8;
m14_mem[8'h15] <= 8'hd6;
m14_mem[8'h16] <= 8'hc4;
m14_mem[8'h17] <= 8'hca;
m14_mem[8'h18] <= 8'h90;
m14_mem[8'h19] <= 8'h9e;
m14_mem[8'h1a] <= 8'h8c;
m14_mem[8'h1b] <= 8'h82;
m14_mem[8'h1c] <= 8'ha8;
m14_mem[8'h1d] <= 8'ha6;
m14_mem[8'h1e] <= 8'hb4;
m14_mem[8'h1f] <= 8'hba;
m14_mem[8'h20] <= 8'hdb;
m14_mem[8'h21] <= 8'hd5;
m14_mem[8'h22] <= 8'hc7;
m14_mem[8'h23] <= 8'hc9;
m14_mem[8'h24] <= 8'he3;
m14_mem[8'h25] <= 8'hed;
m14_mem[8'h26] <= 8'hff;
m14_mem[8'h27] <= 8'hf1;
m14_mem[8'h28] <= 8'hab;
m14_mem[8'h29] <= 8'ha5;
m14_mem[8'h2a] <= 8'hb7;
m14_mem[8'h2b] <= 8'hb9;
m14_mem[8'h2c] <= 8'h93;
m14_mem[8'h2d] <= 8'h9d;
m14_mem[8'h2e] <= 8'h8f;
m14_mem[8'h2f] <= 8'h81;
m14_mem[8'h30] <= 8'h3b;
m14_mem[8'h31] <= 8'h35;
m14_mem[8'h32] <= 8'h27;
m14_mem[8'h33] <= 8'h29;
m14_mem[8'h34] <= 8'h03;
m14_mem[8'h35] <= 8'h0d;
m14_mem[8'h36] <= 8'h1f;
m14_mem[8'h37] <= 8'h11;
m14_mem[8'h38] <= 8'h4b;
m14_mem[8'h39] <= 8'h45;
m14_mem[8'h3a] <= 8'h57;
m14_mem[8'h3b] <= 8'h59;
m14_mem[8'h3c] <= 8'h73;
m14_mem[8'h3d] <= 8'h7d;
m14_mem[8'h3e] <= 8'h6f;
m14_mem[8'h3f] <= 8'h61;
m14_mem[8'h40] <= 8'had;
m14_mem[8'h41] <= 8'ha3;
m14_mem[8'h42] <= 8'hb1;
m14_mem[8'h43] <= 8'hbf;
m14_mem[8'h44] <= 8'h95;
m14_mem[8'h45] <= 8'h9b;
m14_mem[8'h46] <= 8'h89;
m14_mem[8'h47] <= 8'h87;
m14_mem[8'h48] <= 8'hdd;
m14_mem[8'h49] <= 8'hd3;
m14_mem[8'h4a] <= 8'hc1;
m14_mem[8'h4b] <= 8'hcf;
m14_mem[8'h4c] <= 8'he5;
m14_mem[8'h4d] <= 8'heb;
m14_mem[8'h4e] <= 8'hf9;
m14_mem[8'h4f] <= 8'hf7;
m14_mem[8'h50] <= 8'h4d;
m14_mem[8'h51] <= 8'h43;
m14_mem[8'h52] <= 8'h51;
m14_mem[8'h53] <= 8'h5f;
m14_mem[8'h54] <= 8'h75;
m14_mem[8'h55] <= 8'h7b;
m14_mem[8'h56] <= 8'h69;
m14_mem[8'h57] <= 8'h67;
m14_mem[8'h58] <= 8'h3d;
m14_mem[8'h59] <= 8'h33;
m14_mem[8'h5a] <= 8'h21;
m14_mem[8'h5b] <= 8'h2f;
m14_mem[8'h5c] <= 8'h05;
m14_mem[8'h5d] <= 8'h0b;
m14_mem[8'h5e] <= 8'h19;
m14_mem[8'h5f] <= 8'h17;
m14_mem[8'h60] <= 8'h76;
m14_mem[8'h61] <= 8'h78;
m14_mem[8'h62] <= 8'h6a;
m14_mem[8'h63] <= 8'h64;
m14_mem[8'h64] <= 8'h4e;
m14_mem[8'h65] <= 8'h40;
m14_mem[8'h66] <= 8'h52;
m14_mem[8'h67] <= 8'h5c;
m14_mem[8'h68] <= 8'h06;
m14_mem[8'h69] <= 8'h08;
m14_mem[8'h6a] <= 8'h1a;
m14_mem[8'h6b] <= 8'h14;
m14_mem[8'h6c] <= 8'h3e;
m14_mem[8'h6d] <= 8'h30;
m14_mem[8'h6e] <= 8'h22;
m14_mem[8'h6f] <= 8'h2c;
m14_mem[8'h70] <= 8'h96;
m14_mem[8'h71] <= 8'h98;
m14_mem[8'h72] <= 8'h8a;
m14_mem[8'h73] <= 8'h84;
m14_mem[8'h74] <= 8'hae;
m14_mem[8'h75] <= 8'ha0;
m14_mem[8'h76] <= 8'hb2;
m14_mem[8'h77] <= 8'hbc;
m14_mem[8'h78] <= 8'he6;
m14_mem[8'h79] <= 8'he8;
m14_mem[8'h7a] <= 8'hfa;
m14_mem[8'h7b] <= 8'hf4;
m14_mem[8'h7c] <= 8'hde;
m14_mem[8'h7d] <= 8'hd0;
m14_mem[8'h7e] <= 8'hc2;
m14_mem[8'h7f] <= 8'hcc;
m14_mem[8'h80] <= 8'h41;
m14_mem[8'h81] <= 8'h4f;
m14_mem[8'h82] <= 8'h5d;
m14_mem[8'h83] <= 8'h53;
m14_mem[8'h84] <= 8'h79;
m14_mem[8'h85] <= 8'h77;
m14_mem[8'h86] <= 8'h65;
m14_mem[8'h87] <= 8'h6b;
m14_mem[8'h88] <= 8'h31;
m14_mem[8'h89] <= 8'h3f;
m14_mem[8'h8a] <= 8'h2d;
m14_mem[8'h8b] <= 8'h23;
m14_mem[8'h8c] <= 8'h09;
m14_mem[8'h8d] <= 8'h07;
m14_mem[8'h8e] <= 8'h15;
m14_mem[8'h8f] <= 8'h1b;
m14_mem[8'h90] <= 8'ha1;
m14_mem[8'h91] <= 8'haf;
m14_mem[8'h92] <= 8'hbd;
m14_mem[8'h93] <= 8'hb3;
m14_mem[8'h94] <= 8'h99;
m14_mem[8'h95] <= 8'h97;
m14_mem[8'h96] <= 8'h85;
m14_mem[8'h97] <= 8'h8b;
m14_mem[8'h98] <= 8'hd1;
m14_mem[8'h99] <= 8'hdf;
m14_mem[8'h9a] <= 8'hcd;
m14_mem[8'h9b] <= 8'hc3;
m14_mem[8'h9c] <= 8'he9;
m14_mem[8'h9d] <= 8'he7;
m14_mem[8'h9e] <= 8'hf5;
m14_mem[8'h9f] <= 8'hfb;
m14_mem[8'ha0] <= 8'h9a;
m14_mem[8'ha1] <= 8'h94;
m14_mem[8'ha2] <= 8'h86;
m14_mem[8'ha3] <= 8'h88;
m14_mem[8'ha4] <= 8'ha2;
m14_mem[8'ha5] <= 8'hac;
m14_mem[8'ha6] <= 8'hbe;
m14_mem[8'ha7] <= 8'hb0;
m14_mem[8'ha8] <= 8'hea;
m14_mem[8'ha9] <= 8'he4;
m14_mem[8'haa] <= 8'hf6;
m14_mem[8'hab] <= 8'hf8;
m14_mem[8'hac] <= 8'hd2;
m14_mem[8'had] <= 8'hdc;
m14_mem[8'hae] <= 8'hce;
m14_mem[8'haf] <= 8'hc0;
m14_mem[8'hb0] <= 8'h7a;
m14_mem[8'hb1] <= 8'h74;
m14_mem[8'hb2] <= 8'h66;
m14_mem[8'hb3] <= 8'h68;
m14_mem[8'hb4] <= 8'h42;
m14_mem[8'hb5] <= 8'h4c;
m14_mem[8'hb6] <= 8'h5e;
m14_mem[8'hb7] <= 8'h50;
m14_mem[8'hb8] <= 8'h0a;
m14_mem[8'hb9] <= 8'h04;
m14_mem[8'hba] <= 8'h16;
m14_mem[8'hbb] <= 8'h18;
m14_mem[8'hbc] <= 8'h32;
m14_mem[8'hbd] <= 8'h3c;
m14_mem[8'hbe] <= 8'h2e;
m14_mem[8'hbf] <= 8'h20;
m14_mem[8'hc0] <= 8'hec;
m14_mem[8'hc1] <= 8'he2;
m14_mem[8'hc2] <= 8'hf0;
m14_mem[8'hc3] <= 8'hfe;
m14_mem[8'hc4] <= 8'hd4;
m14_mem[8'hc5] <= 8'hda;
m14_mem[8'hc6] <= 8'hc8;
m14_mem[8'hc7] <= 8'hc6;
m14_mem[8'hc8] <= 8'h9c;
m14_mem[8'hc9] <= 8'h92;
m14_mem[8'hca] <= 8'h80;
m14_mem[8'hcb] <= 8'h8e;
m14_mem[8'hcc] <= 8'ha4;
m14_mem[8'hcd] <= 8'haa;
m14_mem[8'hce] <= 8'hb8;
m14_mem[8'hcf] <= 8'hb6;
m14_mem[8'hd0] <= 8'h0c;
m14_mem[8'hd1] <= 8'h02;
m14_mem[8'hd2] <= 8'h10;
m14_mem[8'hd3] <= 8'h1e;
m14_mem[8'hd4] <= 8'h34;
m14_mem[8'hd5] <= 8'h3a;
m14_mem[8'hd6] <= 8'h28;
m14_mem[8'hd7] <= 8'h26;
m14_mem[8'hd8] <= 8'h7c;
m14_mem[8'hd9] <= 8'h72;
m14_mem[8'hda] <= 8'h60;
m14_mem[8'hdb] <= 8'h6e;
m14_mem[8'hdc] <= 8'h44;
m14_mem[8'hdd] <= 8'h4a;
m14_mem[8'hde] <= 8'h58;
m14_mem[8'hdf] <= 8'h56;
m14_mem[8'he0] <= 8'h37;
m14_mem[8'he1] <= 8'h39;
m14_mem[8'he2] <= 8'h2b;
m14_mem[8'he3] <= 8'h25;
m14_mem[8'he4] <= 8'h0f;
m14_mem[8'he5] <= 8'h01;
m14_mem[8'he6] <= 8'h13;
m14_mem[8'he7] <= 8'h1d;
m14_mem[8'he8] <= 8'h47;
m14_mem[8'he9] <= 8'h49;
m14_mem[8'hea] <= 8'h5b;
m14_mem[8'heb] <= 8'h55;
m14_mem[8'hec] <= 8'h7f;
m14_mem[8'hed] <= 8'h71;
m14_mem[8'hee] <= 8'h63;
m14_mem[8'hef] <= 8'h6d;
m14_mem[8'hf0] <= 8'hd7;
m14_mem[8'hf1] <= 8'hd9;
m14_mem[8'hf2] <= 8'hcb;
m14_mem[8'hf3] <= 8'hc5;
m14_mem[8'hf4] <= 8'hef;
m14_mem[8'hf5] <= 8'he1;
m14_mem[8'hf6] <= 8'hf3;
m14_mem[8'hf7] <= 8'hfd;
m14_mem[8'hf8] <= 8'ha7;
m14_mem[8'hf9] <= 8'ha9;
m14_mem[8'hfa] <= 8'hbb;
m14_mem[8'hfb] <= 8'hb5;
m14_mem[8'hfc] <= 8'h9f;
m14_mem[8'hfd] <= 8'h91;
m14_mem[8'hfe] <= 8'h83;
m14_mem[8'hff] <= 8'h8d;
end  


endmodule
